// Verilog netlist produced by program LSE :  version Diamond (64-bit) 3.12.0.240.2
// Netlist written on Thu Aug 17 18:53:52 2023
//
// Verilog Description of module RingOscillatorGenerate
//

module RingOscillatorGenerate (en, run, out3, out5, out7, out101, 
            out1001, out4999, out1000, out1001_M) /* synthesis syn_module_defined=1 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(61[8:30])
    input en;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(63[9:11])
    output run;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(64[10:13])
    output out3;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(65[10:14])
    output out5;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(65[16:20])
    output out7;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(65[22:26])
    output out101;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(65[28:34])
    output out1001;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(65[36:43])
    output out4999;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(65[45:52])
    output out1000;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(65[54:61])
    output out1001_M;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(65[63:72])
    
    wire out3_c /* synthesis alspreserve=1 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(65[10:14])
    
    wire run_c_c, n229, VCC_net, GND_net;
    
    VHI i60 (.Z(VCC_net));
    OB out1000_pad (.I(GND_net), .O(out1000));   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(65[54:61])
    TSALL TSALL_INST (.TSALL(GND_net));
    \RingOscillatorModule(N=1001)  ring1001_M (.run_c_c(run_c_c), .n229(n229)) /* synthesis syn_module_defined=1 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(78[35:60])
    PUR PUR_INST (.PUR(VCC_net));
    defparam PUR_INST.RST_PULSE = 1;
    VLO i4 (.Z(GND_net));
    OB out4999_pad (.I(GND_net), .O(out4999));   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(65[45:52])
    OB out1001_pad (.I(GND_net), .O(out1001));   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(65[36:43])
    GSR GSR_INST (.GSR(VCC_net));
    OB out101_pad (.I(GND_net), .O(out101));   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(65[28:34])
    OB out7_pad (.I(GND_net), .O(out7));   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(65[22:26])
    IB run_c_pad (.I(en), .O(run_c_c));   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(63[9:11])
    OB out5_pad (.I(GND_net), .O(out5));   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(65[16:20])
    OB out3_pad (.I(out3_c), .O(out3));   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(65[10:14])
    OB run_pad (.I(run_c_c), .O(run));   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(64[10:13])
    OB out1001_M_pad (.I(n229), .O(out1001_M));   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(65[63:72])
    \RingOscillatorBase(N=3)  ring3 (.out3_c(out3_c), .run_c_c(run_c_c)) /* synthesis syn_module_defined=1 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(72[30:45])
    
endmodule
//
// Verilog Description of module TSALL
// module not written out since it is a black-box. 
//

//
// Verilog Description of module \RingOscillatorModule(N=1001) 
//

module \RingOscillatorModule(N=1001)  (run_c_c, n229) /* synthesis syn_module_defined=1 */ ;
    input run_c_c;
    output n229;
    
    wire notGate_0 /* synthesis alspreserve=1 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(25[15:22])
    wire notGate_1000 /* synthesis alspreserve=1 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(25[15:22])
    wire notGate_999 /* synthesis alspreserve=1 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(25[15:22])
    wire notGate_998 /* synthesis alspreserve=1 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(25[15:22])
    wire notGate_997 /* synthesis alspreserve=1 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(25[15:22])
    wire notGate_996 /* synthesis alspreserve=1 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(25[15:22])
    wire notGate_995 /* synthesis alspreserve=1 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(25[15:22])
    wire notGate_994 /* synthesis alspreserve=1 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(25[15:22])
    wire notGate_993 /* synthesis alspreserve=1 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(25[15:22])
    wire notGate_992 /* synthesis alspreserve=1 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(25[15:22])
    wire notGate_991 /* synthesis alspreserve=1 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(25[15:22])
    wire notGate_990 /* synthesis alspreserve=1 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(25[15:22])
    wire notGate_989 /* synthesis alspreserve=1 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(25[15:22])
    wire notGate_988 /* synthesis alspreserve=1 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(25[15:22])
    wire notGate_987 /* synthesis alspreserve=1 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(25[15:22])
    wire notGate_986 /* synthesis alspreserve=1 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(25[15:22])
    wire notGate_985 /* synthesis alspreserve=1 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(25[15:22])
    wire notGate_984 /* synthesis alspreserve=1 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(25[15:22])
    wire notGate_983 /* synthesis alspreserve=1 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(25[15:22])
    wire notGate_982 /* synthesis alspreserve=1 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(25[15:22])
    wire notGate_981 /* synthesis alspreserve=1 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(25[15:22])
    wire notGate_980 /* synthesis alspreserve=1 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(25[15:22])
    wire notGate_979 /* synthesis alspreserve=1 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(25[15:22])
    wire notGate_978 /* synthesis alspreserve=1 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(25[15:22])
    wire notGate_977 /* synthesis alspreserve=1 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(25[15:22])
    wire notGate_976 /* synthesis alspreserve=1 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(25[15:22])
    wire notGate_975 /* synthesis alspreserve=1 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(25[15:22])
    wire notGate_974 /* synthesis alspreserve=1 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(25[15:22])
    wire notGate_973 /* synthesis alspreserve=1 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(25[15:22])
    wire notGate_972 /* synthesis alspreserve=1 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(25[15:22])
    wire notGate_971 /* synthesis alspreserve=1 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(25[15:22])
    wire notGate_970 /* synthesis alspreserve=1 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(25[15:22])
    wire notGate_969 /* synthesis alspreserve=1 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(25[15:22])
    wire notGate_968 /* synthesis alspreserve=1 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(25[15:22])
    wire notGate_967 /* synthesis alspreserve=1 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(25[15:22])
    wire notGate_966 /* synthesis alspreserve=1 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(25[15:22])
    wire notGate_965 /* synthesis alspreserve=1 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(25[15:22])
    wire notGate_964 /* synthesis alspreserve=1 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(25[15:22])
    wire notGate_963 /* synthesis alspreserve=1 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(25[15:22])
    wire notGate_962 /* synthesis alspreserve=1 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(25[15:22])
    wire notGate_961 /* synthesis alspreserve=1 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(25[15:22])
    wire notGate_960 /* synthesis alspreserve=1 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(25[15:22])
    wire notGate_959 /* synthesis alspreserve=1 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(25[15:22])
    wire notGate_958 /* synthesis alspreserve=1 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(25[15:22])
    wire notGate_957 /* synthesis alspreserve=1 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(25[15:22])
    wire notGate_956 /* synthesis alspreserve=1 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(25[15:22])
    wire notGate_955 /* synthesis alspreserve=1 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(25[15:22])
    wire notGate_954 /* synthesis alspreserve=1 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(25[15:22])
    wire notGate_953 /* synthesis alspreserve=1 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(25[15:22])
    wire notGate_952 /* synthesis alspreserve=1 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(25[15:22])
    wire notGate_951 /* synthesis alspreserve=1 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(25[15:22])
    wire notGate_950 /* synthesis alspreserve=1 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(25[15:22])
    wire notGate_949 /* synthesis alspreserve=1 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(25[15:22])
    wire notGate_948 /* synthesis alspreserve=1 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(25[15:22])
    wire notGate_947 /* synthesis alspreserve=1 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(25[15:22])
    wire notGate_946 /* synthesis alspreserve=1 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(25[15:22])
    wire notGate_945 /* synthesis alspreserve=1 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(25[15:22])
    wire notGate_944 /* synthesis alspreserve=1 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(25[15:22])
    wire notGate_943 /* synthesis alspreserve=1 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(25[15:22])
    wire notGate_942 /* synthesis alspreserve=1 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(25[15:22])
    wire notGate_941 /* synthesis alspreserve=1 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(25[15:22])
    wire notGate_940 /* synthesis alspreserve=1 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(25[15:22])
    wire notGate_939 /* synthesis alspreserve=1 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(25[15:22])
    wire notGate_938 /* synthesis alspreserve=1 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(25[15:22])
    wire notGate_937 /* synthesis alspreserve=1 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(25[15:22])
    wire notGate_936 /* synthesis alspreserve=1 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(25[15:22])
    wire notGate_935 /* synthesis alspreserve=1 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(25[15:22])
    wire notGate_934 /* synthesis alspreserve=1 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(25[15:22])
    wire notGate_933 /* synthesis alspreserve=1 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(25[15:22])
    wire notGate_932 /* synthesis alspreserve=1 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(25[15:22])
    wire notGate_931 /* synthesis alspreserve=1 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(25[15:22])
    wire notGate_930 /* synthesis alspreserve=1 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(25[15:22])
    wire notGate_929 /* synthesis alspreserve=1 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(25[15:22])
    wire notGate_928 /* synthesis alspreserve=1 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(25[15:22])
    wire notGate_927 /* synthesis alspreserve=1 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(25[15:22])
    wire notGate_926 /* synthesis alspreserve=1 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(25[15:22])
    wire notGate_925 /* synthesis alspreserve=1 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(25[15:22])
    wire notGate_924 /* synthesis alspreserve=1 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(25[15:22])
    wire notGate_923 /* synthesis alspreserve=1 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(25[15:22])
    wire notGate_922 /* synthesis alspreserve=1 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(25[15:22])
    wire notGate_921 /* synthesis alspreserve=1 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(25[15:22])
    wire notGate_920 /* synthesis alspreserve=1 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(25[15:22])
    wire notGate_919 /* synthesis alspreserve=1 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(25[15:22])
    wire notGate_918 /* synthesis alspreserve=1 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(25[15:22])
    wire notGate_917 /* synthesis alspreserve=1 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(25[15:22])
    wire notGate_916 /* synthesis alspreserve=1 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(25[15:22])
    wire notGate_915 /* synthesis alspreserve=1 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(25[15:22])
    wire notGate_914 /* synthesis alspreserve=1 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(25[15:22])
    wire notGate_913 /* synthesis alspreserve=1 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(25[15:22])
    wire notGate_912 /* synthesis alspreserve=1 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(25[15:22])
    wire notGate_911 /* synthesis alspreserve=1 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(25[15:22])
    wire notGate_910 /* synthesis alspreserve=1 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(25[15:22])
    wire notGate_909 /* synthesis alspreserve=1 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(25[15:22])
    wire notGate_908 /* synthesis alspreserve=1 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(25[15:22])
    wire notGate_907 /* synthesis alspreserve=1 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(25[15:22])
    wire notGate_906 /* synthesis alspreserve=1 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(25[15:22])
    wire notGate_905 /* synthesis alspreserve=1 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(25[15:22])
    wire notGate_904 /* synthesis alspreserve=1 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(25[15:22])
    wire notGate_903 /* synthesis alspreserve=1 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(25[15:22])
    wire notGate_902 /* synthesis alspreserve=1 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(25[15:22])
    wire notGate_901 /* synthesis alspreserve=1 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(25[15:22])
    wire notGate_900 /* synthesis alspreserve=1 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(25[15:22])
    wire notGate_899 /* synthesis alspreserve=1 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(25[15:22])
    wire notGate_898 /* synthesis alspreserve=1 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(25[15:22])
    wire notGate_897 /* synthesis alspreserve=1 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(25[15:22])
    wire notGate_896 /* synthesis alspreserve=1 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(25[15:22])
    wire notGate_895 /* synthesis alspreserve=1 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(25[15:22])
    wire notGate_894 /* synthesis alspreserve=1 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(25[15:22])
    wire notGate_893 /* synthesis alspreserve=1 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(25[15:22])
    wire notGate_892 /* synthesis alspreserve=1 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(25[15:22])
    wire notGate_891 /* synthesis alspreserve=1 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(25[15:22])
    wire notGate_890 /* synthesis alspreserve=1 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(25[15:22])
    wire notGate_889 /* synthesis alspreserve=1 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(25[15:22])
    wire notGate_888 /* synthesis alspreserve=1 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(25[15:22])
    wire notGate_887 /* synthesis alspreserve=1 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(25[15:22])
    wire notGate_886 /* synthesis alspreserve=1 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(25[15:22])
    wire notGate_885 /* synthesis alspreserve=1 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(25[15:22])
    wire notGate_884 /* synthesis alspreserve=1 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(25[15:22])
    wire notGate_883 /* synthesis alspreserve=1 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(25[15:22])
    wire notGate_882 /* synthesis alspreserve=1 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(25[15:22])
    wire notGate_881 /* synthesis alspreserve=1 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(25[15:22])
    wire notGate_880 /* synthesis alspreserve=1 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(25[15:22])
    wire notGate_879 /* synthesis alspreserve=1 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(25[15:22])
    wire notGate_878 /* synthesis alspreserve=1 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(25[15:22])
    wire notGate_877 /* synthesis alspreserve=1 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(25[15:22])
    wire notGate_876 /* synthesis alspreserve=1 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(25[15:22])
    wire notGate_875 /* synthesis alspreserve=1 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(25[15:22])
    wire notGate_874 /* synthesis alspreserve=1 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(25[15:22])
    wire notGate_873 /* synthesis alspreserve=1 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(25[15:22])
    wire notGate_872 /* synthesis alspreserve=1 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(25[15:22])
    wire notGate_871 /* synthesis alspreserve=1 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(25[15:22])
    wire notGate_870 /* synthesis alspreserve=1 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(25[15:22])
    wire notGate_869 /* synthesis alspreserve=1 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(25[15:22])
    wire notGate_868 /* synthesis alspreserve=1 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(25[15:22])
    wire notGate_867 /* synthesis alspreserve=1 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(25[15:22])
    wire notGate_866 /* synthesis alspreserve=1 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(25[15:22])
    wire notGate_865 /* synthesis alspreserve=1 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(25[15:22])
    wire notGate_864 /* synthesis alspreserve=1 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(25[15:22])
    wire notGate_863 /* synthesis alspreserve=1 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(25[15:22])
    wire notGate_862 /* synthesis alspreserve=1 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(25[15:22])
    wire notGate_861 /* synthesis alspreserve=1 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(25[15:22])
    wire notGate_860 /* synthesis alspreserve=1 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(25[15:22])
    wire notGate_859 /* synthesis alspreserve=1 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(25[15:22])
    wire notGate_858 /* synthesis alspreserve=1 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(25[15:22])
    wire notGate_857 /* synthesis alspreserve=1 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(25[15:22])
    wire notGate_856 /* synthesis alspreserve=1 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(25[15:22])
    wire notGate_855 /* synthesis alspreserve=1 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(25[15:22])
    wire notGate_854 /* synthesis alspreserve=1 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(25[15:22])
    wire notGate_853 /* synthesis alspreserve=1 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(25[15:22])
    wire notGate_852 /* synthesis alspreserve=1 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(25[15:22])
    wire notGate_851 /* synthesis alspreserve=1 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(25[15:22])
    wire notGate_850 /* synthesis alspreserve=1 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(25[15:22])
    wire notGate_849 /* synthesis alspreserve=1 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(25[15:22])
    wire notGate_848 /* synthesis alspreserve=1 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(25[15:22])
    wire notGate_847 /* synthesis alspreserve=1 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(25[15:22])
    wire notGate_846 /* synthesis alspreserve=1 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(25[15:22])
    wire notGate_845 /* synthesis alspreserve=1 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(25[15:22])
    wire notGate_844 /* synthesis alspreserve=1 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(25[15:22])
    wire notGate_843 /* synthesis alspreserve=1 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(25[15:22])
    wire notGate_842 /* synthesis alspreserve=1 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(25[15:22])
    wire notGate_841 /* synthesis alspreserve=1 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(25[15:22])
    wire notGate_840 /* synthesis alspreserve=1 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(25[15:22])
    wire notGate_839 /* synthesis alspreserve=1 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(25[15:22])
    wire notGate_838 /* synthesis alspreserve=1 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(25[15:22])
    wire notGate_837 /* synthesis alspreserve=1 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(25[15:22])
    wire notGate_836 /* synthesis alspreserve=1 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(25[15:22])
    wire notGate_835 /* synthesis alspreserve=1 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(25[15:22])
    wire notGate_834 /* synthesis alspreserve=1 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(25[15:22])
    wire notGate_833 /* synthesis alspreserve=1 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(25[15:22])
    wire notGate_832 /* synthesis alspreserve=1 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(25[15:22])
    wire notGate_831 /* synthesis alspreserve=1 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(25[15:22])
    wire notGate_830 /* synthesis alspreserve=1 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(25[15:22])
    wire notGate_829 /* synthesis alspreserve=1 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(25[15:22])
    wire notGate_828 /* synthesis alspreserve=1 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(25[15:22])
    wire notGate_827 /* synthesis alspreserve=1 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(25[15:22])
    wire notGate_826 /* synthesis alspreserve=1 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(25[15:22])
    wire notGate_825 /* synthesis alspreserve=1 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(25[15:22])
    wire notGate_824 /* synthesis alspreserve=1 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(25[15:22])
    wire notGate_823 /* synthesis alspreserve=1 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(25[15:22])
    wire notGate_822 /* synthesis alspreserve=1 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(25[15:22])
    wire notGate_821 /* synthesis alspreserve=1 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(25[15:22])
    wire notGate_820 /* synthesis alspreserve=1 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(25[15:22])
    wire notGate_819 /* synthesis alspreserve=1 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(25[15:22])
    wire notGate_818 /* synthesis alspreserve=1 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(25[15:22])
    wire notGate_817 /* synthesis alspreserve=1 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(25[15:22])
    wire notGate_816 /* synthesis alspreserve=1 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(25[15:22])
    wire notGate_815 /* synthesis alspreserve=1 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(25[15:22])
    wire notGate_814 /* synthesis alspreserve=1 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(25[15:22])
    wire notGate_813 /* synthesis alspreserve=1 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(25[15:22])
    wire notGate_812 /* synthesis alspreserve=1 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(25[15:22])
    wire notGate_811 /* synthesis alspreserve=1 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(25[15:22])
    wire notGate_810 /* synthesis alspreserve=1 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(25[15:22])
    wire notGate_809 /* synthesis alspreserve=1 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(25[15:22])
    wire notGate_808 /* synthesis alspreserve=1 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(25[15:22])
    wire notGate_807 /* synthesis alspreserve=1 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(25[15:22])
    wire notGate_806 /* synthesis alspreserve=1 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(25[15:22])
    wire notGate_805 /* synthesis alspreserve=1 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(25[15:22])
    wire notGate_804 /* synthesis alspreserve=1 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(25[15:22])
    wire notGate_803 /* synthesis alspreserve=1 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(25[15:22])
    wire notGate_802 /* synthesis alspreserve=1 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(25[15:22])
    wire notGate_801 /* synthesis alspreserve=1 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(25[15:22])
    wire notGate_800 /* synthesis alspreserve=1 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(25[15:22])
    wire notGate_799 /* synthesis alspreserve=1 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(25[15:22])
    wire notGate_798 /* synthesis alspreserve=1 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(25[15:22])
    wire notGate_797 /* synthesis alspreserve=1 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(25[15:22])
    wire notGate_796 /* synthesis alspreserve=1 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(25[15:22])
    wire notGate_795 /* synthesis alspreserve=1 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(25[15:22])
    wire notGate_794 /* synthesis alspreserve=1 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(25[15:22])
    wire notGate_793 /* synthesis alspreserve=1 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(25[15:22])
    wire notGate_792 /* synthesis alspreserve=1 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(25[15:22])
    wire notGate_791 /* synthesis alspreserve=1 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(25[15:22])
    wire notGate_790 /* synthesis alspreserve=1 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(25[15:22])
    wire notGate_789 /* synthesis alspreserve=1 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(25[15:22])
    wire notGate_788 /* synthesis alspreserve=1 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(25[15:22])
    wire notGate_787 /* synthesis alspreserve=1 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(25[15:22])
    wire notGate_786 /* synthesis alspreserve=1 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(25[15:22])
    wire notGate_785 /* synthesis alspreserve=1 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(25[15:22])
    wire notGate_784 /* synthesis alspreserve=1 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(25[15:22])
    wire notGate_783 /* synthesis alspreserve=1 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(25[15:22])
    wire notGate_782 /* synthesis alspreserve=1 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(25[15:22])
    wire notGate_781 /* synthesis alspreserve=1 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(25[15:22])
    wire notGate_780 /* synthesis alspreserve=1 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(25[15:22])
    wire notGate_779 /* synthesis alspreserve=1 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(25[15:22])
    wire notGate_778 /* synthesis alspreserve=1 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(25[15:22])
    wire notGate_777 /* synthesis alspreserve=1 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(25[15:22])
    wire notGate_776 /* synthesis alspreserve=1 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(25[15:22])
    wire notGate_775 /* synthesis alspreserve=1 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(25[15:22])
    wire notGate_774 /* synthesis alspreserve=1 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(25[15:22])
    wire notGate_773 /* synthesis alspreserve=1 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(25[15:22])
    wire notGate_772 /* synthesis alspreserve=1 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(25[15:22])
    wire notGate_771 /* synthesis alspreserve=1 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(25[15:22])
    wire notGate_770 /* synthesis alspreserve=1 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(25[15:22])
    wire notGate_769 /* synthesis alspreserve=1 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(25[15:22])
    wire notGate_768 /* synthesis alspreserve=1 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(25[15:22])
    wire notGate_767 /* synthesis alspreserve=1 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(25[15:22])
    wire notGate_766 /* synthesis alspreserve=1 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(25[15:22])
    wire notGate_765 /* synthesis alspreserve=1 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(25[15:22])
    wire notGate_764 /* synthesis alspreserve=1 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(25[15:22])
    wire notGate_763 /* synthesis alspreserve=1 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(25[15:22])
    wire notGate_762 /* synthesis alspreserve=1 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(25[15:22])
    wire notGate_761 /* synthesis alspreserve=1 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(25[15:22])
    wire notGate_760 /* synthesis alspreserve=1 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(25[15:22])
    wire notGate_759 /* synthesis alspreserve=1 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(25[15:22])
    wire notGate_758 /* synthesis alspreserve=1 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(25[15:22])
    wire notGate_757 /* synthesis alspreserve=1 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(25[15:22])
    wire notGate_756 /* synthesis alspreserve=1 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(25[15:22])
    wire notGate_755 /* synthesis alspreserve=1 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(25[15:22])
    wire notGate_754 /* synthesis alspreserve=1 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(25[15:22])
    wire notGate_753 /* synthesis alspreserve=1 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(25[15:22])
    wire notGate_752 /* synthesis alspreserve=1 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(25[15:22])
    wire notGate_751 /* synthesis alspreserve=1 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(25[15:22])
    wire notGate_750 /* synthesis alspreserve=1 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(25[15:22])
    wire notGate_749 /* synthesis alspreserve=1 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(25[15:22])
    wire notGate_748 /* synthesis alspreserve=1 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(25[15:22])
    wire notGate_747 /* synthesis alspreserve=1 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(25[15:22])
    wire notGate_746 /* synthesis alspreserve=1 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(25[15:22])
    wire notGate_745 /* synthesis alspreserve=1 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(25[15:22])
    wire notGate_744 /* synthesis alspreserve=1 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(25[15:22])
    wire notGate_743 /* synthesis alspreserve=1 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(25[15:22])
    wire notGate_742 /* synthesis alspreserve=1 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(25[15:22])
    wire notGate_741 /* synthesis alspreserve=1 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(25[15:22])
    wire notGate_740 /* synthesis alspreserve=1 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(25[15:22])
    wire notGate_739 /* synthesis alspreserve=1 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(25[15:22])
    wire notGate_738 /* synthesis alspreserve=1 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(25[15:22])
    wire notGate_737 /* synthesis alspreserve=1 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(25[15:22])
    wire notGate_736 /* synthesis alspreserve=1 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(25[15:22])
    wire notGate_735 /* synthesis alspreserve=1 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(25[15:22])
    wire notGate_734 /* synthesis alspreserve=1 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(25[15:22])
    wire notGate_733 /* synthesis alspreserve=1 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(25[15:22])
    wire notGate_732 /* synthesis alspreserve=1 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(25[15:22])
    wire notGate_731 /* synthesis alspreserve=1 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(25[15:22])
    wire notGate_730 /* synthesis alspreserve=1 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(25[15:22])
    wire notGate_729 /* synthesis alspreserve=1 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(25[15:22])
    wire notGate_728 /* synthesis alspreserve=1 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(25[15:22])
    wire notGate_727 /* synthesis alspreserve=1 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(25[15:22])
    wire notGate_726 /* synthesis alspreserve=1 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(25[15:22])
    wire notGate_725 /* synthesis alspreserve=1 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(25[15:22])
    wire notGate_724 /* synthesis alspreserve=1 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(25[15:22])
    wire notGate_723 /* synthesis alspreserve=1 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(25[15:22])
    wire notGate_722 /* synthesis alspreserve=1 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(25[15:22])
    wire notGate_721 /* synthesis alspreserve=1 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(25[15:22])
    wire notGate_720 /* synthesis alspreserve=1 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(25[15:22])
    wire notGate_719 /* synthesis alspreserve=1 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(25[15:22])
    wire notGate_718 /* synthesis alspreserve=1 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(25[15:22])
    wire notGate_717 /* synthesis alspreserve=1 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(25[15:22])
    wire notGate_716 /* synthesis alspreserve=1 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(25[15:22])
    wire notGate_715 /* synthesis alspreserve=1 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(25[15:22])
    wire notGate_714 /* synthesis alspreserve=1 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(25[15:22])
    wire notGate_713 /* synthesis alspreserve=1 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(25[15:22])
    wire notGate_712 /* synthesis alspreserve=1 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(25[15:22])
    wire notGate_711 /* synthesis alspreserve=1 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(25[15:22])
    wire notGate_710 /* synthesis alspreserve=1 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(25[15:22])
    wire notGate_709 /* synthesis alspreserve=1 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(25[15:22])
    wire notGate_708 /* synthesis alspreserve=1 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(25[15:22])
    wire notGate_707 /* synthesis alspreserve=1 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(25[15:22])
    wire notGate_706 /* synthesis alspreserve=1 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(25[15:22])
    wire notGate_705 /* synthesis alspreserve=1 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(25[15:22])
    wire notGate_704 /* synthesis alspreserve=1 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(25[15:22])
    wire notGate_703 /* synthesis alspreserve=1 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(25[15:22])
    wire notGate_702 /* synthesis alspreserve=1 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(25[15:22])
    wire notGate_701 /* synthesis alspreserve=1 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(25[15:22])
    wire notGate_700 /* synthesis alspreserve=1 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(25[15:22])
    wire notGate_699 /* synthesis alspreserve=1 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(25[15:22])
    wire notGate_698 /* synthesis alspreserve=1 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(25[15:22])
    wire notGate_697 /* synthesis alspreserve=1 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(25[15:22])
    wire notGate_696 /* synthesis alspreserve=1 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(25[15:22])
    wire notGate_695 /* synthesis alspreserve=1 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(25[15:22])
    wire notGate_694 /* synthesis alspreserve=1 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(25[15:22])
    wire notGate_693 /* synthesis alspreserve=1 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(25[15:22])
    wire notGate_692 /* synthesis alspreserve=1 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(25[15:22])
    wire notGate_691 /* synthesis alspreserve=1 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(25[15:22])
    wire notGate_690 /* synthesis alspreserve=1 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(25[15:22])
    wire notGate_689 /* synthesis alspreserve=1 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(25[15:22])
    wire notGate_688 /* synthesis alspreserve=1 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(25[15:22])
    wire notGate_687 /* synthesis alspreserve=1 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(25[15:22])
    wire notGate_686 /* synthesis alspreserve=1 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(25[15:22])
    wire notGate_685 /* synthesis alspreserve=1 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(25[15:22])
    wire notGate_684 /* synthesis alspreserve=1 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(25[15:22])
    wire notGate_683 /* synthesis alspreserve=1 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(25[15:22])
    wire notGate_682 /* synthesis alspreserve=1 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(25[15:22])
    wire notGate_681 /* synthesis alspreserve=1 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(25[15:22])
    wire notGate_680 /* synthesis alspreserve=1 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(25[15:22])
    wire notGate_679 /* synthesis alspreserve=1 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(25[15:22])
    wire notGate_678 /* synthesis alspreserve=1 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(25[15:22])
    wire notGate_677 /* synthesis alspreserve=1 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(25[15:22])
    wire notGate_676 /* synthesis alspreserve=1 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(25[15:22])
    wire notGate_675 /* synthesis alspreserve=1 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(25[15:22])
    wire notGate_674 /* synthesis alspreserve=1 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(25[15:22])
    wire notGate_673 /* synthesis alspreserve=1 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(25[15:22])
    wire notGate_672 /* synthesis alspreserve=1 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(25[15:22])
    wire notGate_671 /* synthesis alspreserve=1 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(25[15:22])
    wire notGate_670 /* synthesis alspreserve=1 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(25[15:22])
    wire notGate_669 /* synthesis alspreserve=1 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(25[15:22])
    wire notGate_668 /* synthesis alspreserve=1 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(25[15:22])
    wire notGate_667 /* synthesis alspreserve=1 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(25[15:22])
    wire notGate_666 /* synthesis alspreserve=1 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(25[15:22])
    wire notGate_665 /* synthesis alspreserve=1 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(25[15:22])
    wire notGate_664 /* synthesis alspreserve=1 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(25[15:22])
    wire notGate_663 /* synthesis alspreserve=1 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(25[15:22])
    wire notGate_662 /* synthesis alspreserve=1 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(25[15:22])
    wire notGate_661 /* synthesis alspreserve=1 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(25[15:22])
    wire notGate_660 /* synthesis alspreserve=1 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(25[15:22])
    wire notGate_659 /* synthesis alspreserve=1 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(25[15:22])
    wire notGate_658 /* synthesis alspreserve=1 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(25[15:22])
    wire notGate_657 /* synthesis alspreserve=1 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(25[15:22])
    wire notGate_656 /* synthesis alspreserve=1 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(25[15:22])
    wire notGate_655 /* synthesis alspreserve=1 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(25[15:22])
    wire notGate_654 /* synthesis alspreserve=1 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(25[15:22])
    wire notGate_653 /* synthesis alspreserve=1 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(25[15:22])
    wire notGate_652 /* synthesis alspreserve=1 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(25[15:22])
    wire notGate_651 /* synthesis alspreserve=1 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(25[15:22])
    wire notGate_650 /* synthesis alspreserve=1 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(25[15:22])
    wire notGate_649 /* synthesis alspreserve=1 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(25[15:22])
    wire notGate_648 /* synthesis alspreserve=1 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(25[15:22])
    wire notGate_647 /* synthesis alspreserve=1 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(25[15:22])
    wire notGate_646 /* synthesis alspreserve=1 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(25[15:22])
    wire notGate_645 /* synthesis alspreserve=1 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(25[15:22])
    wire notGate_644 /* synthesis alspreserve=1 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(25[15:22])
    wire notGate_643 /* synthesis alspreserve=1 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(25[15:22])
    wire notGate_642 /* synthesis alspreserve=1 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(25[15:22])
    wire notGate_641 /* synthesis alspreserve=1 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(25[15:22])
    wire notGate_640 /* synthesis alspreserve=1 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(25[15:22])
    wire notGate_639 /* synthesis alspreserve=1 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(25[15:22])
    wire notGate_638 /* synthesis alspreserve=1 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(25[15:22])
    wire notGate_637 /* synthesis alspreserve=1 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(25[15:22])
    wire notGate_636 /* synthesis alspreserve=1 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(25[15:22])
    wire notGate_635 /* synthesis alspreserve=1 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(25[15:22])
    wire notGate_634 /* synthesis alspreserve=1 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(25[15:22])
    wire notGate_633 /* synthesis alspreserve=1 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(25[15:22])
    wire notGate_632 /* synthesis alspreserve=1 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(25[15:22])
    wire notGate_631 /* synthesis alspreserve=1 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(25[15:22])
    wire notGate_630 /* synthesis alspreserve=1 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(25[15:22])
    wire notGate_629 /* synthesis alspreserve=1 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(25[15:22])
    wire notGate_628 /* synthesis alspreserve=1 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(25[15:22])
    wire notGate_627 /* synthesis alspreserve=1 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(25[15:22])
    wire notGate_626 /* synthesis alspreserve=1 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(25[15:22])
    wire notGate_625 /* synthesis alspreserve=1 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(25[15:22])
    wire notGate_624 /* synthesis alspreserve=1 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(25[15:22])
    wire notGate_623 /* synthesis alspreserve=1 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(25[15:22])
    wire notGate_622 /* synthesis alspreserve=1 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(25[15:22])
    wire notGate_621 /* synthesis alspreserve=1 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(25[15:22])
    wire notGate_620 /* synthesis alspreserve=1 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(25[15:22])
    wire notGate_619 /* synthesis alspreserve=1 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(25[15:22])
    wire notGate_618 /* synthesis alspreserve=1 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(25[15:22])
    wire notGate_617 /* synthesis alspreserve=1 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(25[15:22])
    wire notGate_616 /* synthesis alspreserve=1 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(25[15:22])
    wire notGate_615 /* synthesis alspreserve=1 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(25[15:22])
    wire notGate_614 /* synthesis alspreserve=1 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(25[15:22])
    wire notGate_613 /* synthesis alspreserve=1 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(25[15:22])
    wire notGate_612 /* synthesis alspreserve=1 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(25[15:22])
    wire notGate_611 /* synthesis alspreserve=1 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(25[15:22])
    wire notGate_610 /* synthesis alspreserve=1 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(25[15:22])
    wire notGate_609 /* synthesis alspreserve=1 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(25[15:22])
    wire notGate_608 /* synthesis alspreserve=1 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(25[15:22])
    wire notGate_607 /* synthesis alspreserve=1 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(25[15:22])
    wire notGate_606 /* synthesis alspreserve=1 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(25[15:22])
    wire notGate_605 /* synthesis alspreserve=1 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(25[15:22])
    wire notGate_604 /* synthesis alspreserve=1 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(25[15:22])
    wire notGate_603 /* synthesis alspreserve=1 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(25[15:22])
    wire notGate_602 /* synthesis alspreserve=1 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(25[15:22])
    wire notGate_601 /* synthesis alspreserve=1 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(25[15:22])
    wire notGate_600 /* synthesis alspreserve=1 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(25[15:22])
    wire notGate_599 /* synthesis alspreserve=1 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(25[15:22])
    wire notGate_598 /* synthesis alspreserve=1 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(25[15:22])
    wire notGate_597 /* synthesis alspreserve=1 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(25[15:22])
    wire notGate_596 /* synthesis alspreserve=1 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(25[15:22])
    wire notGate_595 /* synthesis alspreserve=1 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(25[15:22])
    wire notGate_594 /* synthesis alspreserve=1 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(25[15:22])
    wire notGate_593 /* synthesis alspreserve=1 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(25[15:22])
    wire notGate_592 /* synthesis alspreserve=1 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(25[15:22])
    wire notGate_591 /* synthesis alspreserve=1 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(25[15:22])
    wire notGate_590 /* synthesis alspreserve=1 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(25[15:22])
    wire notGate_589 /* synthesis alspreserve=1 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(25[15:22])
    wire notGate_588 /* synthesis alspreserve=1 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(25[15:22])
    wire notGate_587 /* synthesis alspreserve=1 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(25[15:22])
    wire notGate_586 /* synthesis alspreserve=1 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(25[15:22])
    wire notGate_585 /* synthesis alspreserve=1 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(25[15:22])
    wire notGate_584 /* synthesis alspreserve=1 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(25[15:22])
    wire notGate_583 /* synthesis alspreserve=1 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(25[15:22])
    wire notGate_582 /* synthesis alspreserve=1 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(25[15:22])
    wire notGate_581 /* synthesis alspreserve=1 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(25[15:22])
    wire notGate_580 /* synthesis alspreserve=1 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(25[15:22])
    wire notGate_579 /* synthesis alspreserve=1 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(25[15:22])
    wire notGate_578 /* synthesis alspreserve=1 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(25[15:22])
    wire notGate_577 /* synthesis alspreserve=1 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(25[15:22])
    wire notGate_576 /* synthesis alspreserve=1 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(25[15:22])
    wire notGate_575 /* synthesis alspreserve=1 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(25[15:22])
    wire notGate_574 /* synthesis alspreserve=1 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(25[15:22])
    wire notGate_573 /* synthesis alspreserve=1 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(25[15:22])
    wire notGate_572 /* synthesis alspreserve=1 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(25[15:22])
    wire notGate_571 /* synthesis alspreserve=1 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(25[15:22])
    wire notGate_570 /* synthesis alspreserve=1 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(25[15:22])
    wire notGate_569 /* synthesis alspreserve=1 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(25[15:22])
    wire notGate_568 /* synthesis alspreserve=1 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(25[15:22])
    wire notGate_567 /* synthesis alspreserve=1 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(25[15:22])
    wire notGate_566 /* synthesis alspreserve=1 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(25[15:22])
    wire notGate_565 /* synthesis alspreserve=1 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(25[15:22])
    wire notGate_564 /* synthesis alspreserve=1 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(25[15:22])
    wire notGate_563 /* synthesis alspreserve=1 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(25[15:22])
    wire notGate_562 /* synthesis alspreserve=1 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(25[15:22])
    wire notGate_561 /* synthesis alspreserve=1 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(25[15:22])
    wire notGate_560 /* synthesis alspreserve=1 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(25[15:22])
    wire notGate_559 /* synthesis alspreserve=1 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(25[15:22])
    wire notGate_558 /* synthesis alspreserve=1 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(25[15:22])
    wire notGate_557 /* synthesis alspreserve=1 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(25[15:22])
    wire notGate_556 /* synthesis alspreserve=1 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(25[15:22])
    wire notGate_555 /* synthesis alspreserve=1 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(25[15:22])
    wire notGate_554 /* synthesis alspreserve=1 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(25[15:22])
    wire notGate_553 /* synthesis alspreserve=1 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(25[15:22])
    wire notGate_552 /* synthesis alspreserve=1 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(25[15:22])
    wire notGate_551 /* synthesis alspreserve=1 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(25[15:22])
    wire notGate_550 /* synthesis alspreserve=1 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(25[15:22])
    wire notGate_549 /* synthesis alspreserve=1 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(25[15:22])
    wire notGate_548 /* synthesis alspreserve=1 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(25[15:22])
    wire notGate_547 /* synthesis alspreserve=1 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(25[15:22])
    wire notGate_546 /* synthesis alspreserve=1 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(25[15:22])
    wire notGate_545 /* synthesis alspreserve=1 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(25[15:22])
    wire notGate_544 /* synthesis alspreserve=1 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(25[15:22])
    wire notGate_543 /* synthesis alspreserve=1 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(25[15:22])
    wire notGate_542 /* synthesis alspreserve=1 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(25[15:22])
    wire notGate_541 /* synthesis alspreserve=1 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(25[15:22])
    wire notGate_540 /* synthesis alspreserve=1 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(25[15:22])
    wire notGate_539 /* synthesis alspreserve=1 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(25[15:22])
    wire notGate_538 /* synthesis alspreserve=1 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(25[15:22])
    wire notGate_537 /* synthesis alspreserve=1 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(25[15:22])
    wire notGate_536 /* synthesis alspreserve=1 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(25[15:22])
    wire notGate_535 /* synthesis alspreserve=1 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(25[15:22])
    wire notGate_534 /* synthesis alspreserve=1 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(25[15:22])
    wire notGate_533 /* synthesis alspreserve=1 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(25[15:22])
    wire notGate_532 /* synthesis alspreserve=1 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(25[15:22])
    wire notGate_531 /* synthesis alspreserve=1 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(25[15:22])
    wire notGate_530 /* synthesis alspreserve=1 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(25[15:22])
    wire notGate_529 /* synthesis alspreserve=1 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(25[15:22])
    wire notGate_528 /* synthesis alspreserve=1 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(25[15:22])
    wire notGate_527 /* synthesis alspreserve=1 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(25[15:22])
    wire notGate_526 /* synthesis alspreserve=1 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(25[15:22])
    wire notGate_525 /* synthesis alspreserve=1 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(25[15:22])
    wire notGate_524 /* synthesis alspreserve=1 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(25[15:22])
    wire notGate_523 /* synthesis alspreserve=1 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(25[15:22])
    wire notGate_522 /* synthesis alspreserve=1 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(25[15:22])
    wire notGate_521 /* synthesis alspreserve=1 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(25[15:22])
    wire notGate_520 /* synthesis alspreserve=1 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(25[15:22])
    wire notGate_519 /* synthesis alspreserve=1 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(25[15:22])
    wire notGate_518 /* synthesis alspreserve=1 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(25[15:22])
    wire notGate_517 /* synthesis alspreserve=1 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(25[15:22])
    wire notGate_516 /* synthesis alspreserve=1 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(25[15:22])
    wire notGate_515 /* synthesis alspreserve=1 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(25[15:22])
    wire notGate_514 /* synthesis alspreserve=1 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(25[15:22])
    wire notGate_513 /* synthesis alspreserve=1 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(25[15:22])
    wire notGate_512 /* synthesis alspreserve=1 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(25[15:22])
    wire notGate_511 /* synthesis alspreserve=1 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(25[15:22])
    wire notGate_510 /* synthesis alspreserve=1 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(25[15:22])
    wire notGate_509 /* synthesis alspreserve=1 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(25[15:22])
    wire notGate_508 /* synthesis alspreserve=1 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(25[15:22])
    wire notGate_507 /* synthesis alspreserve=1 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(25[15:22])
    wire notGate_506 /* synthesis alspreserve=1 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(25[15:22])
    wire notGate_505 /* synthesis alspreserve=1 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(25[15:22])
    wire notGate_504 /* synthesis alspreserve=1 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(25[15:22])
    wire notGate_503 /* synthesis alspreserve=1 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(25[15:22])
    wire notGate_502 /* synthesis alspreserve=1 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(25[15:22])
    wire notGate_501 /* synthesis alspreserve=1 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(25[15:22])
    wire notGate_500 /* synthesis alspreserve=1 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(25[15:22])
    wire notGate_499 /* synthesis alspreserve=1 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(25[15:22])
    wire notGate_498 /* synthesis alspreserve=1 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(25[15:22])
    wire notGate_497 /* synthesis alspreserve=1 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(25[15:22])
    wire notGate_496 /* synthesis alspreserve=1 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(25[15:22])
    wire notGate_495 /* synthesis alspreserve=1 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(25[15:22])
    wire notGate_494 /* synthesis alspreserve=1 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(25[15:22])
    wire notGate_493 /* synthesis alspreserve=1 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(25[15:22])
    wire notGate_492 /* synthesis alspreserve=1 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(25[15:22])
    wire notGate_491 /* synthesis alspreserve=1 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(25[15:22])
    wire notGate_490 /* synthesis alspreserve=1 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(25[15:22])
    wire notGate_489 /* synthesis alspreserve=1 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(25[15:22])
    wire notGate_488 /* synthesis alspreserve=1 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(25[15:22])
    wire notGate_487 /* synthesis alspreserve=1 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(25[15:22])
    wire notGate_486 /* synthesis alspreserve=1 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(25[15:22])
    wire notGate_485 /* synthesis alspreserve=1 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(25[15:22])
    wire notGate_484 /* synthesis alspreserve=1 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(25[15:22])
    wire notGate_483 /* synthesis alspreserve=1 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(25[15:22])
    wire notGate_482 /* synthesis alspreserve=1 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(25[15:22])
    wire notGate_481 /* synthesis alspreserve=1 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(25[15:22])
    wire notGate_480 /* synthesis alspreserve=1 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(25[15:22])
    wire notGate_479 /* synthesis alspreserve=1 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(25[15:22])
    wire notGate_478 /* synthesis alspreserve=1 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(25[15:22])
    wire notGate_477 /* synthesis alspreserve=1 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(25[15:22])
    wire notGate_476 /* synthesis alspreserve=1 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(25[15:22])
    wire notGate_475 /* synthesis alspreserve=1 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(25[15:22])
    wire notGate_474 /* synthesis alspreserve=1 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(25[15:22])
    wire notGate_473 /* synthesis alspreserve=1 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(25[15:22])
    wire notGate_472 /* synthesis alspreserve=1 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(25[15:22])
    wire notGate_471 /* synthesis alspreserve=1 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(25[15:22])
    wire notGate_470 /* synthesis alspreserve=1 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(25[15:22])
    wire notGate_469 /* synthesis alspreserve=1 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(25[15:22])
    wire notGate_468 /* synthesis alspreserve=1 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(25[15:22])
    wire notGate_467 /* synthesis alspreserve=1 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(25[15:22])
    wire notGate_466 /* synthesis alspreserve=1 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(25[15:22])
    wire notGate_465 /* synthesis alspreserve=1 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(25[15:22])
    wire notGate_464 /* synthesis alspreserve=1 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(25[15:22])
    wire notGate_463 /* synthesis alspreserve=1 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(25[15:22])
    wire notGate_462 /* synthesis alspreserve=1 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(25[15:22])
    wire notGate_461 /* synthesis alspreserve=1 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(25[15:22])
    wire notGate_460 /* synthesis alspreserve=1 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(25[15:22])
    wire notGate_459 /* synthesis alspreserve=1 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(25[15:22])
    wire notGate_458 /* synthesis alspreserve=1 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(25[15:22])
    wire notGate_457 /* synthesis alspreserve=1 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(25[15:22])
    wire notGate_456 /* synthesis alspreserve=1 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(25[15:22])
    wire notGate_455 /* synthesis alspreserve=1 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(25[15:22])
    wire notGate_454 /* synthesis alspreserve=1 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(25[15:22])
    wire notGate_453 /* synthesis alspreserve=1 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(25[15:22])
    wire notGate_452 /* synthesis alspreserve=1 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(25[15:22])
    wire notGate_451 /* synthesis alspreserve=1 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(25[15:22])
    wire notGate_450 /* synthesis alspreserve=1 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(25[15:22])
    wire notGate_449 /* synthesis alspreserve=1 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(25[15:22])
    wire notGate_448 /* synthesis alspreserve=1 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(25[15:22])
    wire notGate_447 /* synthesis alspreserve=1 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(25[15:22])
    wire notGate_446 /* synthesis alspreserve=1 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(25[15:22])
    wire notGate_445 /* synthesis alspreserve=1 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(25[15:22])
    wire notGate_444 /* synthesis alspreserve=1 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(25[15:22])
    wire notGate_443 /* synthesis alspreserve=1 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(25[15:22])
    wire notGate_442 /* synthesis alspreserve=1 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(25[15:22])
    wire notGate_441 /* synthesis alspreserve=1 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(25[15:22])
    wire notGate_440 /* synthesis alspreserve=1 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(25[15:22])
    wire notGate_439 /* synthesis alspreserve=1 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(25[15:22])
    wire notGate_438 /* synthesis alspreserve=1 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(25[15:22])
    wire notGate_437 /* synthesis alspreserve=1 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(25[15:22])
    wire notGate_436 /* synthesis alspreserve=1 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(25[15:22])
    wire notGate_435 /* synthesis alspreserve=1 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(25[15:22])
    wire notGate_434 /* synthesis alspreserve=1 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(25[15:22])
    wire notGate_433 /* synthesis alspreserve=1 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(25[15:22])
    wire notGate_432 /* synthesis alspreserve=1 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(25[15:22])
    wire notGate_431 /* synthesis alspreserve=1 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(25[15:22])
    wire notGate_430 /* synthesis alspreserve=1 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(25[15:22])
    wire notGate_429 /* synthesis alspreserve=1 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(25[15:22])
    wire notGate_428 /* synthesis alspreserve=1 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(25[15:22])
    wire notGate_427 /* synthesis alspreserve=1 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(25[15:22])
    wire notGate_426 /* synthesis alspreserve=1 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(25[15:22])
    wire notGate_425 /* synthesis alspreserve=1 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(25[15:22])
    wire notGate_424 /* synthesis alspreserve=1 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(25[15:22])
    wire notGate_423 /* synthesis alspreserve=1 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(25[15:22])
    wire notGate_422 /* synthesis alspreserve=1 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(25[15:22])
    wire notGate_421 /* synthesis alspreserve=1 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(25[15:22])
    wire notGate_420 /* synthesis alspreserve=1 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(25[15:22])
    wire notGate_419 /* synthesis alspreserve=1 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(25[15:22])
    wire notGate_418 /* synthesis alspreserve=1 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(25[15:22])
    wire notGate_417 /* synthesis alspreserve=1 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(25[15:22])
    wire notGate_416 /* synthesis alspreserve=1 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(25[15:22])
    wire notGate_415 /* synthesis alspreserve=1 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(25[15:22])
    wire notGate_414 /* synthesis alspreserve=1 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(25[15:22])
    wire notGate_413 /* synthesis alspreserve=1 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(25[15:22])
    wire notGate_412 /* synthesis alspreserve=1 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(25[15:22])
    wire notGate_411 /* synthesis alspreserve=1 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(25[15:22])
    wire notGate_410 /* synthesis alspreserve=1 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(25[15:22])
    wire notGate_409 /* synthesis alspreserve=1 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(25[15:22])
    wire notGate_408 /* synthesis alspreserve=1 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(25[15:22])
    wire notGate_407 /* synthesis alspreserve=1 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(25[15:22])
    wire notGate_406 /* synthesis alspreserve=1 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(25[15:22])
    wire notGate_405 /* synthesis alspreserve=1 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(25[15:22])
    wire notGate_404 /* synthesis alspreserve=1 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(25[15:22])
    wire notGate_403 /* synthesis alspreserve=1 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(25[15:22])
    wire notGate_402 /* synthesis alspreserve=1 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(25[15:22])
    wire notGate_401 /* synthesis alspreserve=1 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(25[15:22])
    wire notGate_400 /* synthesis alspreserve=1 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(25[15:22])
    wire notGate_399 /* synthesis alspreserve=1 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(25[15:22])
    wire notGate_398 /* synthesis alspreserve=1 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(25[15:22])
    wire notGate_397 /* synthesis alspreserve=1 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(25[15:22])
    wire notGate_396 /* synthesis alspreserve=1 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(25[15:22])
    wire notGate_395 /* synthesis alspreserve=1 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(25[15:22])
    wire notGate_394 /* synthesis alspreserve=1 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(25[15:22])
    wire notGate_393 /* synthesis alspreserve=1 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(25[15:22])
    wire notGate_392 /* synthesis alspreserve=1 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(25[15:22])
    wire notGate_391 /* synthesis alspreserve=1 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(25[15:22])
    wire notGate_390 /* synthesis alspreserve=1 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(25[15:22])
    wire notGate_389 /* synthesis alspreserve=1 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(25[15:22])
    wire notGate_388 /* synthesis alspreserve=1 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(25[15:22])
    wire notGate_387 /* synthesis alspreserve=1 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(25[15:22])
    wire notGate_386 /* synthesis alspreserve=1 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(25[15:22])
    wire notGate_385 /* synthesis alspreserve=1 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(25[15:22])
    wire notGate_384 /* synthesis alspreserve=1 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(25[15:22])
    wire notGate_383 /* synthesis alspreserve=1 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(25[15:22])
    wire notGate_382 /* synthesis alspreserve=1 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(25[15:22])
    wire notGate_381 /* synthesis alspreserve=1 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(25[15:22])
    wire notGate_380 /* synthesis alspreserve=1 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(25[15:22])
    wire notGate_379 /* synthesis alspreserve=1 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(25[15:22])
    wire notGate_378 /* synthesis alspreserve=1 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(25[15:22])
    wire notGate_377 /* synthesis alspreserve=1 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(25[15:22])
    wire notGate_376 /* synthesis alspreserve=1 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(25[15:22])
    wire notGate_375 /* synthesis alspreserve=1 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(25[15:22])
    wire notGate_374 /* synthesis alspreserve=1 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(25[15:22])
    wire notGate_373 /* synthesis alspreserve=1 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(25[15:22])
    wire notGate_372 /* synthesis alspreserve=1 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(25[15:22])
    wire notGate_371 /* synthesis alspreserve=1 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(25[15:22])
    wire notGate_370 /* synthesis alspreserve=1 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(25[15:22])
    wire notGate_369 /* synthesis alspreserve=1 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(25[15:22])
    wire notGate_368 /* synthesis alspreserve=1 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(25[15:22])
    wire notGate_367 /* synthesis alspreserve=1 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(25[15:22])
    wire notGate_366 /* synthesis alspreserve=1 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(25[15:22])
    wire notGate_365 /* synthesis alspreserve=1 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(25[15:22])
    wire notGate_364 /* synthesis alspreserve=1 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(25[15:22])
    wire notGate_363 /* synthesis alspreserve=1 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(25[15:22])
    wire notGate_362 /* synthesis alspreserve=1 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(25[15:22])
    wire notGate_361 /* synthesis alspreserve=1 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(25[15:22])
    wire notGate_360 /* synthesis alspreserve=1 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(25[15:22])
    wire notGate_359 /* synthesis alspreserve=1 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(25[15:22])
    wire notGate_358 /* synthesis alspreserve=1 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(25[15:22])
    wire notGate_357 /* synthesis alspreserve=1 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(25[15:22])
    wire notGate_356 /* synthesis alspreserve=1 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(25[15:22])
    wire notGate_355 /* synthesis alspreserve=1 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(25[15:22])
    wire notGate_354 /* synthesis alspreserve=1 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(25[15:22])
    wire notGate_353 /* synthesis alspreserve=1 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(25[15:22])
    wire notGate_352 /* synthesis alspreserve=1 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(25[15:22])
    wire notGate_351 /* synthesis alspreserve=1 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(25[15:22])
    wire notGate_350 /* synthesis alspreserve=1 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(25[15:22])
    wire notGate_349 /* synthesis alspreserve=1 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(25[15:22])
    wire notGate_348 /* synthesis alspreserve=1 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(25[15:22])
    wire notGate_347 /* synthesis alspreserve=1 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(25[15:22])
    wire notGate_346 /* synthesis alspreserve=1 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(25[15:22])
    wire notGate_345 /* synthesis alspreserve=1 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(25[15:22])
    wire notGate_344 /* synthesis alspreserve=1 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(25[15:22])
    wire notGate_343 /* synthesis alspreserve=1 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(25[15:22])
    wire notGate_342 /* synthesis alspreserve=1 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(25[15:22])
    wire notGate_341 /* synthesis alspreserve=1 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(25[15:22])
    wire notGate_340 /* synthesis alspreserve=1 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(25[15:22])
    wire notGate_339 /* synthesis alspreserve=1 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(25[15:22])
    wire notGate_338 /* synthesis alspreserve=1 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(25[15:22])
    wire notGate_337 /* synthesis alspreserve=1 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(25[15:22])
    wire notGate_336 /* synthesis alspreserve=1 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(25[15:22])
    wire notGate_335 /* synthesis alspreserve=1 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(25[15:22])
    wire notGate_334 /* synthesis alspreserve=1 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(25[15:22])
    wire notGate_333 /* synthesis alspreserve=1 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(25[15:22])
    wire notGate_332 /* synthesis alspreserve=1 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(25[15:22])
    wire notGate_331 /* synthesis alspreserve=1 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(25[15:22])
    wire notGate_330 /* synthesis alspreserve=1 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(25[15:22])
    wire notGate_329 /* synthesis alspreserve=1 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(25[15:22])
    wire notGate_328 /* synthesis alspreserve=1 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(25[15:22])
    wire notGate_327 /* synthesis alspreserve=1 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(25[15:22])
    wire notGate_326 /* synthesis alspreserve=1 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(25[15:22])
    wire notGate_325 /* synthesis alspreserve=1 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(25[15:22])
    wire notGate_324 /* synthesis alspreserve=1 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(25[15:22])
    wire notGate_323 /* synthesis alspreserve=1 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(25[15:22])
    wire notGate_322 /* synthesis alspreserve=1 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(25[15:22])
    wire notGate_321 /* synthesis alspreserve=1 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(25[15:22])
    wire notGate_320 /* synthesis alspreserve=1 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(25[15:22])
    wire notGate_319 /* synthesis alspreserve=1 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(25[15:22])
    wire notGate_318 /* synthesis alspreserve=1 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(25[15:22])
    wire notGate_317 /* synthesis alspreserve=1 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(25[15:22])
    wire notGate_316 /* synthesis alspreserve=1 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(25[15:22])
    wire notGate_315 /* synthesis alspreserve=1 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(25[15:22])
    wire notGate_314 /* synthesis alspreserve=1 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(25[15:22])
    wire notGate_313 /* synthesis alspreserve=1 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(25[15:22])
    wire notGate_312 /* synthesis alspreserve=1 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(25[15:22])
    wire notGate_311 /* synthesis alspreserve=1 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(25[15:22])
    wire notGate_310 /* synthesis alspreserve=1 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(25[15:22])
    wire notGate_309 /* synthesis alspreserve=1 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(25[15:22])
    wire notGate_308 /* synthesis alspreserve=1 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(25[15:22])
    wire notGate_307 /* synthesis alspreserve=1 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(25[15:22])
    wire notGate_306 /* synthesis alspreserve=1 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(25[15:22])
    wire notGate_305 /* synthesis alspreserve=1 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(25[15:22])
    wire notGate_304 /* synthesis alspreserve=1 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(25[15:22])
    wire notGate_303 /* synthesis alspreserve=1 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(25[15:22])
    wire notGate_302 /* synthesis alspreserve=1 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(25[15:22])
    wire notGate_301 /* synthesis alspreserve=1 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(25[15:22])
    wire notGate_300 /* synthesis alspreserve=1 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(25[15:22])
    wire notGate_299 /* synthesis alspreserve=1 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(25[15:22])
    wire notGate_298 /* synthesis alspreserve=1 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(25[15:22])
    wire notGate_297 /* synthesis alspreserve=1 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(25[15:22])
    wire notGate_296 /* synthesis alspreserve=1 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(25[15:22])
    wire notGate_295 /* synthesis alspreserve=1 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(25[15:22])
    wire notGate_294 /* synthesis alspreserve=1 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(25[15:22])
    wire notGate_293 /* synthesis alspreserve=1 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(25[15:22])
    wire notGate_292 /* synthesis alspreserve=1 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(25[15:22])
    wire notGate_291 /* synthesis alspreserve=1 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(25[15:22])
    wire notGate_290 /* synthesis alspreserve=1 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(25[15:22])
    wire notGate_289 /* synthesis alspreserve=1 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(25[15:22])
    wire notGate_288 /* synthesis alspreserve=1 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(25[15:22])
    wire notGate_287 /* synthesis alspreserve=1 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(25[15:22])
    wire notGate_286 /* synthesis alspreserve=1 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(25[15:22])
    wire notGate_285 /* synthesis alspreserve=1 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(25[15:22])
    wire notGate_284 /* synthesis alspreserve=1 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(25[15:22])
    wire notGate_283 /* synthesis alspreserve=1 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(25[15:22])
    wire notGate_282 /* synthesis alspreserve=1 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(25[15:22])
    wire notGate_281 /* synthesis alspreserve=1 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(25[15:22])
    wire notGate_280 /* synthesis alspreserve=1 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(25[15:22])
    wire notGate_279 /* synthesis alspreserve=1 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(25[15:22])
    wire notGate_278 /* synthesis alspreserve=1 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(25[15:22])
    wire notGate_277 /* synthesis alspreserve=1 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(25[15:22])
    wire notGate_276 /* synthesis alspreserve=1 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(25[15:22])
    wire notGate_275 /* synthesis alspreserve=1 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(25[15:22])
    wire notGate_274 /* synthesis alspreserve=1 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(25[15:22])
    wire notGate_273 /* synthesis alspreserve=1 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(25[15:22])
    wire notGate_272 /* synthesis alspreserve=1 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(25[15:22])
    wire notGate_271 /* synthesis alspreserve=1 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(25[15:22])
    wire notGate_270 /* synthesis alspreserve=1 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(25[15:22])
    wire notGate_269 /* synthesis alspreserve=1 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(25[15:22])
    wire notGate_268 /* synthesis alspreserve=1 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(25[15:22])
    wire notGate_267 /* synthesis alspreserve=1 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(25[15:22])
    wire notGate_266 /* synthesis alspreserve=1 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(25[15:22])
    wire notGate_265 /* synthesis alspreserve=1 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(25[15:22])
    wire notGate_264 /* synthesis alspreserve=1 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(25[15:22])
    wire notGate_263 /* synthesis alspreserve=1 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(25[15:22])
    wire notGate_262 /* synthesis alspreserve=1 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(25[15:22])
    wire notGate_261 /* synthesis alspreserve=1 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(25[15:22])
    wire notGate_260 /* synthesis alspreserve=1 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(25[15:22])
    wire notGate_259 /* synthesis alspreserve=1 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(25[15:22])
    wire notGate_258 /* synthesis alspreserve=1 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(25[15:22])
    wire notGate_257 /* synthesis alspreserve=1 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(25[15:22])
    wire notGate_256 /* synthesis alspreserve=1 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(25[15:22])
    wire notGate_255 /* synthesis alspreserve=1 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(25[15:22])
    wire notGate_254 /* synthesis alspreserve=1 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(25[15:22])
    wire notGate_253 /* synthesis alspreserve=1 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(25[15:22])
    wire notGate_252 /* synthesis alspreserve=1 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(25[15:22])
    wire notGate_251 /* synthesis alspreserve=1 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(25[15:22])
    wire notGate_250 /* synthesis alspreserve=1 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(25[15:22])
    wire notGate_249 /* synthesis alspreserve=1 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(25[15:22])
    wire notGate_248 /* synthesis alspreserve=1 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(25[15:22])
    wire notGate_247 /* synthesis alspreserve=1 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(25[15:22])
    wire notGate_246 /* synthesis alspreserve=1 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(25[15:22])
    wire notGate_245 /* synthesis alspreserve=1 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(25[15:22])
    wire notGate_244 /* synthesis alspreserve=1 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(25[15:22])
    wire notGate_243 /* synthesis alspreserve=1 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(25[15:22])
    wire notGate_242 /* synthesis alspreserve=1 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(25[15:22])
    wire notGate_241 /* synthesis alspreserve=1 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(25[15:22])
    wire notGate_240 /* synthesis alspreserve=1 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(25[15:22])
    wire notGate_239 /* synthesis alspreserve=1 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(25[15:22])
    wire notGate_238 /* synthesis alspreserve=1 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(25[15:22])
    wire notGate_237 /* synthesis alspreserve=1 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(25[15:22])
    wire notGate_236 /* synthesis alspreserve=1 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(25[15:22])
    wire notGate_235 /* synthesis alspreserve=1 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(25[15:22])
    wire notGate_234 /* synthesis alspreserve=1 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(25[15:22])
    wire notGate_233 /* synthesis alspreserve=1 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(25[15:22])
    wire notGate_232 /* synthesis alspreserve=1 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(25[15:22])
    wire notGate_231 /* synthesis alspreserve=1 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(25[15:22])
    wire notGate_230 /* synthesis alspreserve=1 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(25[15:22])
    wire notGate_229 /* synthesis alspreserve=1 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(25[15:22])
    wire notGate_228 /* synthesis alspreserve=1 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(25[15:22])
    wire notGate_227 /* synthesis alspreserve=1 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(25[15:22])
    wire notGate_226 /* synthesis alspreserve=1 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(25[15:22])
    wire notGate_225 /* synthesis alspreserve=1 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(25[15:22])
    wire notGate_224 /* synthesis alspreserve=1 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(25[15:22])
    wire notGate_223 /* synthesis alspreserve=1 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(25[15:22])
    wire notGate_222 /* synthesis alspreserve=1 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(25[15:22])
    wire notGate_221 /* synthesis alspreserve=1 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(25[15:22])
    wire notGate_220 /* synthesis alspreserve=1 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(25[15:22])
    wire notGate_219 /* synthesis alspreserve=1 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(25[15:22])
    wire notGate_218 /* synthesis alspreserve=1 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(25[15:22])
    wire notGate_217 /* synthesis alspreserve=1 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(25[15:22])
    wire notGate_216 /* synthesis alspreserve=1 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(25[15:22])
    wire notGate_215 /* synthesis alspreserve=1 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(25[15:22])
    wire notGate_214 /* synthesis alspreserve=1 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(25[15:22])
    wire notGate_213 /* synthesis alspreserve=1 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(25[15:22])
    wire notGate_212 /* synthesis alspreserve=1 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(25[15:22])
    wire notGate_211 /* synthesis alspreserve=1 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(25[15:22])
    wire notGate_210 /* synthesis alspreserve=1 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(25[15:22])
    wire notGate_209 /* synthesis alspreserve=1 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(25[15:22])
    wire notGate_208 /* synthesis alspreserve=1 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(25[15:22])
    wire notGate_207 /* synthesis alspreserve=1 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(25[15:22])
    wire notGate_206 /* synthesis alspreserve=1 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(25[15:22])
    wire notGate_205 /* synthesis alspreserve=1 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(25[15:22])
    wire notGate_204 /* synthesis alspreserve=1 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(25[15:22])
    wire notGate_203 /* synthesis alspreserve=1 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(25[15:22])
    wire notGate_202 /* synthesis alspreserve=1 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(25[15:22])
    wire notGate_201 /* synthesis alspreserve=1 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(25[15:22])
    wire notGate_200 /* synthesis alspreserve=1 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(25[15:22])
    wire notGate_199 /* synthesis alspreserve=1 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(25[15:22])
    wire notGate_198 /* synthesis alspreserve=1 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(25[15:22])
    wire notGate_197 /* synthesis alspreserve=1 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(25[15:22])
    wire notGate_196 /* synthesis alspreserve=1 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(25[15:22])
    wire notGate_195 /* synthesis alspreserve=1 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(25[15:22])
    wire notGate_194 /* synthesis alspreserve=1 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(25[15:22])
    wire notGate_193 /* synthesis alspreserve=1 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(25[15:22])
    wire notGate_192 /* synthesis alspreserve=1 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(25[15:22])
    wire notGate_191 /* synthesis alspreserve=1 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(25[15:22])
    wire notGate_190 /* synthesis alspreserve=1 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(25[15:22])
    wire notGate_189 /* synthesis alspreserve=1 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(25[15:22])
    wire notGate_188 /* synthesis alspreserve=1 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(25[15:22])
    wire notGate_187 /* synthesis alspreserve=1 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(25[15:22])
    wire notGate_186 /* synthesis alspreserve=1 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(25[15:22])
    wire notGate_185 /* synthesis alspreserve=1 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(25[15:22])
    wire notGate_184 /* synthesis alspreserve=1 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(25[15:22])
    wire notGate_183 /* synthesis alspreserve=1 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(25[15:22])
    wire notGate_182 /* synthesis alspreserve=1 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(25[15:22])
    wire notGate_181 /* synthesis alspreserve=1 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(25[15:22])
    wire notGate_180 /* synthesis alspreserve=1 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(25[15:22])
    wire notGate_179 /* synthesis alspreserve=1 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(25[15:22])
    wire notGate_178 /* synthesis alspreserve=1 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(25[15:22])
    wire notGate_177 /* synthesis alspreserve=1 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(25[15:22])
    wire notGate_176 /* synthesis alspreserve=1 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(25[15:22])
    wire notGate_175 /* synthesis alspreserve=1 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(25[15:22])
    wire notGate_174 /* synthesis alspreserve=1 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(25[15:22])
    wire notGate_173 /* synthesis alspreserve=1 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(25[15:22])
    wire notGate_172 /* synthesis alspreserve=1 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(25[15:22])
    wire notGate_171 /* synthesis alspreserve=1 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(25[15:22])
    wire notGate_170 /* synthesis alspreserve=1 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(25[15:22])
    wire notGate_169 /* synthesis alspreserve=1 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(25[15:22])
    wire notGate_168 /* synthesis alspreserve=1 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(25[15:22])
    wire notGate_167 /* synthesis alspreserve=1 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(25[15:22])
    wire notGate_166 /* synthesis alspreserve=1 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(25[15:22])
    wire notGate_165 /* synthesis alspreserve=1 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(25[15:22])
    wire notGate_164 /* synthesis alspreserve=1 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(25[15:22])
    wire notGate_163 /* synthesis alspreserve=1 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(25[15:22])
    wire notGate_162 /* synthesis alspreserve=1 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(25[15:22])
    wire notGate_161 /* synthesis alspreserve=1 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(25[15:22])
    wire notGate_160 /* synthesis alspreserve=1 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(25[15:22])
    wire notGate_159 /* synthesis alspreserve=1 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(25[15:22])
    wire notGate_158 /* synthesis alspreserve=1 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(25[15:22])
    wire notGate_157 /* synthesis alspreserve=1 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(25[15:22])
    wire notGate_156 /* synthesis alspreserve=1 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(25[15:22])
    wire notGate_155 /* synthesis alspreserve=1 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(25[15:22])
    wire notGate_154 /* synthesis alspreserve=1 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(25[15:22])
    wire notGate_153 /* synthesis alspreserve=1 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(25[15:22])
    wire notGate_152 /* synthesis alspreserve=1 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(25[15:22])
    wire notGate_151 /* synthesis alspreserve=1 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(25[15:22])
    wire notGate_150 /* synthesis alspreserve=1 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(25[15:22])
    wire notGate_149 /* synthesis alspreserve=1 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(25[15:22])
    wire notGate_148 /* synthesis alspreserve=1 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(25[15:22])
    wire notGate_147 /* synthesis alspreserve=1 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(25[15:22])
    wire notGate_146 /* synthesis alspreserve=1 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(25[15:22])
    wire notGate_145 /* synthesis alspreserve=1 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(25[15:22])
    wire notGate_144 /* synthesis alspreserve=1 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(25[15:22])
    wire notGate_143 /* synthesis alspreserve=1 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(25[15:22])
    wire notGate_142 /* synthesis alspreserve=1 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(25[15:22])
    wire notGate_141 /* synthesis alspreserve=1 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(25[15:22])
    wire notGate_140 /* synthesis alspreserve=1 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(25[15:22])
    wire notGate_139 /* synthesis alspreserve=1 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(25[15:22])
    wire notGate_138 /* synthesis alspreserve=1 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(25[15:22])
    wire notGate_137 /* synthesis alspreserve=1 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(25[15:22])
    wire notGate_136 /* synthesis alspreserve=1 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(25[15:22])
    wire notGate_135 /* synthesis alspreserve=1 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(25[15:22])
    wire notGate_134 /* synthesis alspreserve=1 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(25[15:22])
    wire notGate_133 /* synthesis alspreserve=1 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(25[15:22])
    wire notGate_132 /* synthesis alspreserve=1 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(25[15:22])
    wire notGate_131 /* synthesis alspreserve=1 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(25[15:22])
    wire notGate_130 /* synthesis alspreserve=1 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(25[15:22])
    wire notGate_129 /* synthesis alspreserve=1 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(25[15:22])
    wire notGate_128 /* synthesis alspreserve=1 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(25[15:22])
    wire notGate_127 /* synthesis alspreserve=1 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(25[15:22])
    wire notGate_126 /* synthesis alspreserve=1 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(25[15:22])
    wire notGate_125 /* synthesis alspreserve=1 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(25[15:22])
    wire notGate_124 /* synthesis alspreserve=1 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(25[15:22])
    wire notGate_123 /* synthesis alspreserve=1 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(25[15:22])
    wire notGate_122 /* synthesis alspreserve=1 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(25[15:22])
    wire notGate_121 /* synthesis alspreserve=1 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(25[15:22])
    wire notGate_120 /* synthesis alspreserve=1 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(25[15:22])
    wire notGate_119 /* synthesis alspreserve=1 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(25[15:22])
    wire notGate_118 /* synthesis alspreserve=1 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(25[15:22])
    wire notGate_117 /* synthesis alspreserve=1 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(25[15:22])
    wire notGate_116 /* synthesis alspreserve=1 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(25[15:22])
    wire notGate_115 /* synthesis alspreserve=1 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(25[15:22])
    wire notGate_114 /* synthesis alspreserve=1 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(25[15:22])
    wire notGate_113 /* synthesis alspreserve=1 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(25[15:22])
    wire notGate_112 /* synthesis alspreserve=1 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(25[15:22])
    wire notGate_111 /* synthesis alspreserve=1 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(25[15:22])
    wire notGate_110 /* synthesis alspreserve=1 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(25[15:22])
    wire notGate_109 /* synthesis alspreserve=1 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(25[15:22])
    wire notGate_108 /* synthesis alspreserve=1 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(25[15:22])
    wire notGate_107 /* synthesis alspreserve=1 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(25[15:22])
    wire notGate_106 /* synthesis alspreserve=1 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(25[15:22])
    wire notGate_105 /* synthesis alspreserve=1 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(25[15:22])
    wire notGate_104 /* synthesis alspreserve=1 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(25[15:22])
    wire notGate_103 /* synthesis alspreserve=1 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(25[15:22])
    wire notGate_102 /* synthesis alspreserve=1 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(25[15:22])
    wire notGate_101 /* synthesis alspreserve=1 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(25[15:22])
    wire notGate_100 /* synthesis alspreserve=1 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(25[15:22])
    wire notGate_99 /* synthesis alspreserve=1 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(25[15:22])
    wire notGate_98 /* synthesis alspreserve=1 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(25[15:22])
    wire notGate_97 /* synthesis alspreserve=1 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(25[15:22])
    wire notGate_96 /* synthesis alspreserve=1 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(25[15:22])
    wire notGate_95 /* synthesis alspreserve=1 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(25[15:22])
    wire notGate_94 /* synthesis alspreserve=1 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(25[15:22])
    wire notGate_93 /* synthesis alspreserve=1 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(25[15:22])
    wire notGate_92 /* synthesis alspreserve=1 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(25[15:22])
    wire notGate_91 /* synthesis alspreserve=1 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(25[15:22])
    wire notGate_90 /* synthesis alspreserve=1 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(25[15:22])
    wire notGate_89 /* synthesis alspreserve=1 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(25[15:22])
    wire notGate_88 /* synthesis alspreserve=1 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(25[15:22])
    wire notGate_87 /* synthesis alspreserve=1 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(25[15:22])
    wire notGate_86 /* synthesis alspreserve=1 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(25[15:22])
    wire notGate_85 /* synthesis alspreserve=1 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(25[15:22])
    wire notGate_84 /* synthesis alspreserve=1 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(25[15:22])
    wire notGate_83 /* synthesis alspreserve=1 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(25[15:22])
    wire notGate_82 /* synthesis alspreserve=1 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(25[15:22])
    wire notGate_81 /* synthesis alspreserve=1 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(25[15:22])
    wire notGate_80 /* synthesis alspreserve=1 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(25[15:22])
    wire notGate_79 /* synthesis alspreserve=1 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(25[15:22])
    wire notGate_78 /* synthesis alspreserve=1 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(25[15:22])
    wire notGate_77 /* synthesis alspreserve=1 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(25[15:22])
    wire notGate_76 /* synthesis alspreserve=1 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(25[15:22])
    wire notGate_75 /* synthesis alspreserve=1 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(25[15:22])
    wire notGate_74 /* synthesis alspreserve=1 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(25[15:22])
    wire notGate_73 /* synthesis alspreserve=1 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(25[15:22])
    wire notGate_72 /* synthesis alspreserve=1 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(25[15:22])
    wire notGate_71 /* synthesis alspreserve=1 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(25[15:22])
    wire notGate_70 /* synthesis alspreserve=1 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(25[15:22])
    wire notGate_69 /* synthesis alspreserve=1 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(25[15:22])
    wire notGate_68 /* synthesis alspreserve=1 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(25[15:22])
    wire notGate_67 /* synthesis alspreserve=1 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(25[15:22])
    wire notGate_66 /* synthesis alspreserve=1 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(25[15:22])
    wire notGate_65 /* synthesis alspreserve=1 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(25[15:22])
    wire notGate_64 /* synthesis alspreserve=1 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(25[15:22])
    wire notGate_63 /* synthesis alspreserve=1 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(25[15:22])
    wire notGate_62 /* synthesis alspreserve=1 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(25[15:22])
    wire notGate_61 /* synthesis alspreserve=1 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(25[15:22])
    wire notGate_60 /* synthesis alspreserve=1 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(25[15:22])
    wire notGate_59 /* synthesis alspreserve=1 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(25[15:22])
    wire notGate_58 /* synthesis alspreserve=1 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(25[15:22])
    wire notGate_57 /* synthesis alspreserve=1 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(25[15:22])
    wire notGate_56 /* synthesis alspreserve=1 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(25[15:22])
    wire notGate_55 /* synthesis alspreserve=1 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(25[15:22])
    wire notGate_54 /* synthesis alspreserve=1 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(25[15:22])
    wire notGate_53 /* synthesis alspreserve=1 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(25[15:22])
    wire notGate_52 /* synthesis alspreserve=1 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(25[15:22])
    wire notGate_51 /* synthesis alspreserve=1 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(25[15:22])
    wire notGate_50 /* synthesis alspreserve=1 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(25[15:22])
    wire notGate_49 /* synthesis alspreserve=1 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(25[15:22])
    wire notGate_48 /* synthesis alspreserve=1 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(25[15:22])
    wire notGate_47 /* synthesis alspreserve=1 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(25[15:22])
    wire notGate_46 /* synthesis alspreserve=1 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(25[15:22])
    wire notGate_45 /* synthesis alspreserve=1 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(25[15:22])
    wire notGate_44 /* synthesis alspreserve=1 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(25[15:22])
    wire notGate_43 /* synthesis alspreserve=1 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(25[15:22])
    wire notGate_42 /* synthesis alspreserve=1 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(25[15:22])
    wire notGate_41 /* synthesis alspreserve=1 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(25[15:22])
    wire notGate_40 /* synthesis alspreserve=1 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(25[15:22])
    wire notGate_39 /* synthesis alspreserve=1 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(25[15:22])
    wire notGate_38 /* synthesis alspreserve=1 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(25[15:22])
    wire notGate_37 /* synthesis alspreserve=1 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(25[15:22])
    wire notGate_36 /* synthesis alspreserve=1 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(25[15:22])
    wire notGate_35 /* synthesis alspreserve=1 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(25[15:22])
    wire notGate_34 /* synthesis alspreserve=1 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(25[15:22])
    wire notGate_33 /* synthesis alspreserve=1 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(25[15:22])
    wire notGate_32 /* synthesis alspreserve=1 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(25[15:22])
    wire notGate_31 /* synthesis alspreserve=1 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(25[15:22])
    wire notGate_30 /* synthesis alspreserve=1 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(25[15:22])
    wire notGate_29 /* synthesis alspreserve=1 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(25[15:22])
    wire notGate_28 /* synthesis alspreserve=1 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(25[15:22])
    wire notGate_27 /* synthesis alspreserve=1 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(25[15:22])
    wire notGate_26 /* synthesis alspreserve=1 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(25[15:22])
    wire notGate_25 /* synthesis alspreserve=1 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(25[15:22])
    wire notGate_24 /* synthesis alspreserve=1 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(25[15:22])
    wire notGate_23 /* synthesis alspreserve=1 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(25[15:22])
    wire notGate_22 /* synthesis alspreserve=1 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(25[15:22])
    wire notGate_21 /* synthesis alspreserve=1 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(25[15:22])
    wire notGate_20 /* synthesis alspreserve=1 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(25[15:22])
    wire notGate_19 /* synthesis alspreserve=1 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(25[15:22])
    wire notGate_18 /* synthesis alspreserve=1 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(25[15:22])
    wire notGate_17 /* synthesis alspreserve=1 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(25[15:22])
    wire notGate_16 /* synthesis alspreserve=1 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(25[15:22])
    wire notGate_15 /* synthesis alspreserve=1 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(25[15:22])
    wire notGate_14 /* synthesis alspreserve=1 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(25[15:22])
    wire notGate_13 /* synthesis alspreserve=1 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(25[15:22])
    wire notGate_12 /* synthesis alspreserve=1 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(25[15:22])
    wire notGate_11 /* synthesis alspreserve=1 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(25[15:22])
    wire notGate_10 /* synthesis alspreserve=1 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(25[15:22])
    wire notGate_9 /* synthesis alspreserve=1 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(25[15:22])
    wire notGate_8 /* synthesis alspreserve=1 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(25[15:22])
    wire notGate_7 /* synthesis alspreserve=1 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(25[15:22])
    wire notGate_6 /* synthesis alspreserve=1 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(25[15:22])
    wire notGate_5 /* synthesis alspreserve=1 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(25[15:22])
    wire notGate_4 /* synthesis alspreserve=1 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(25[15:22])
    wire notGate_3 /* synthesis alspreserve=1 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(25[15:22])
    wire notGate_2 /* synthesis alspreserve=1 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(25[15:22])
    wire notGate_1 /* synthesis alspreserve=1 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(25[15:22])
    
    LUT4 en_I_0_2_lut_rep_1 (.A(run_c_c), .B(notGate_1000), .Z(n229)) /* synthesis lut_function=(A (B)) */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(29[18:35])
    defparam en_I_0_2_lut_rep_1.init = 16'h8888;
    LUT4 and_1_I_0_1_lut_2_lut (.A(run_c_c), .B(notGate_1000), .Z(notGate_0)) /* synthesis lut_function=(!(A (B))) */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(29[18:35])
    defparam and_1_I_0_1_lut_2_lut.init = 16'h7777;
    inverter \inverter_chain_9..inv  (.\notGate[8]_keep (notGate_8), .\notGate[9] (notGate_9)) /* synthesis syn_module_defined=1 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(32[13:44])
    inverter_U0 \inverter_chain_99..inv  (.\notGate[98]_keep (notGate_98), 
            .\notGate[99] (notGate_99)) /* synthesis syn_module_defined=1 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(32[13:44])
    inverter_U1 \inverter_chain_999..inv  (.\notGate[998]_keep (notGate_998), 
            .\notGate[999] (notGate_999)) /* synthesis syn_module_defined=1 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(32[13:44])
    inverter_U2 \inverter_chain_998..inv  (.\notGate[997]_keep (notGate_997), 
            .\notGate[998] (notGate_998)) /* synthesis syn_module_defined=1 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(32[13:44])
    inverter_U3 \inverter_chain_997..inv  (.\notGate[996]_keep (notGate_996), 
            .\notGate[997] (notGate_997)) /* synthesis syn_module_defined=1 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(32[13:44])
    inverter_U4 \inverter_chain_996..inv  (.\notGate[995]_keep (notGate_995), 
            .\notGate[996] (notGate_996)) /* synthesis syn_module_defined=1 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(32[13:44])
    inverter_U5 \inverter_chain_995..inv  (.\notGate[994]_keep (notGate_994), 
            .\notGate[995] (notGate_995)) /* synthesis syn_module_defined=1 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(32[13:44])
    inverter_U6 \inverter_chain_994..inv  (.\notGate[993]_keep (notGate_993), 
            .\notGate[994] (notGate_994)) /* synthesis syn_module_defined=1 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(32[13:44])
    inverter_U7 \inverter_chain_993..inv  (.\notGate[992]_keep (notGate_992), 
            .\notGate[993] (notGate_993)) /* synthesis syn_module_defined=1 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(32[13:44])
    inverter_U8 \inverter_chain_992..inv  (.\notGate[991]_keep (notGate_991), 
            .\notGate[992] (notGate_992)) /* synthesis syn_module_defined=1 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(32[13:44])
    inverter_U9 \inverter_chain_991..inv  (.\notGate[990]_keep (notGate_990), 
            .\notGate[991] (notGate_991)) /* synthesis syn_module_defined=1 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(32[13:44])
    inverter_U10 \inverter_chain_990..inv  (.\notGate[989]_keep (notGate_989), 
            .\notGate[990] (notGate_990)) /* synthesis syn_module_defined=1 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(32[13:44])
    inverter_U11 \inverter_chain_98..inv  (.\notGate[97]_keep (notGate_97), 
            .\notGate[98] (notGate_98)) /* synthesis syn_module_defined=1 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(32[13:44])
    inverter_U12 \inverter_chain_989..inv  (.\notGate[988]_keep (notGate_988), 
            .\notGate[989] (notGate_989)) /* synthesis syn_module_defined=1 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(32[13:44])
    inverter_U13 \inverter_chain_988..inv  (.\notGate[987]_keep (notGate_987), 
            .\notGate[988] (notGate_988)) /* synthesis syn_module_defined=1 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(32[13:44])
    inverter_U14 \inverter_chain_987..inv  (.\notGate[986]_keep (notGate_986), 
            .\notGate[987] (notGate_987)) /* synthesis syn_module_defined=1 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(32[13:44])
    inverter_U15 \inverter_chain_986..inv  (.\notGate[985]_keep (notGate_985), 
            .\notGate[986] (notGate_986)) /* synthesis syn_module_defined=1 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(32[13:44])
    inverter_U16 \inverter_chain_985..inv  (.\notGate[984]_keep (notGate_984), 
            .\notGate[985] (notGate_985)) /* synthesis syn_module_defined=1 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(32[13:44])
    inverter_U17 \inverter_chain_984..inv  (.\notGate[983]_keep (notGate_983), 
            .\notGate[984] (notGate_984)) /* synthesis syn_module_defined=1 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(32[13:44])
    inverter_U18 \inverter_chain_983..inv  (.\notGate[982]_keep (notGate_982), 
            .\notGate[983] (notGate_983)) /* synthesis syn_module_defined=1 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(32[13:44])
    inverter_U19 \inverter_chain_982..inv  (.\notGate[981]_keep (notGate_981), 
            .\notGate[982] (notGate_982)) /* synthesis syn_module_defined=1 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(32[13:44])
    inverter_U20 \inverter_chain_981..inv  (.\notGate[980]_keep (notGate_980), 
            .\notGate[981] (notGate_981)) /* synthesis syn_module_defined=1 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(32[13:44])
    inverter_U21 \inverter_chain_980..inv  (.\notGate[979]_keep (notGate_979), 
            .\notGate[980] (notGate_980)) /* synthesis syn_module_defined=1 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(32[13:44])
    inverter_U22 \inverter_chain_97..inv  (.\notGate[96]_keep (notGate_96), 
            .\notGate[97] (notGate_97)) /* synthesis syn_module_defined=1 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(32[13:44])
    inverter_U23 \inverter_chain_979..inv  (.\notGate[978]_keep (notGate_978), 
            .\notGate[979] (notGate_979)) /* synthesis syn_module_defined=1 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(32[13:44])
    inverter_U24 \inverter_chain_978..inv  (.\notGate[977]_keep (notGate_977), 
            .\notGate[978] (notGate_978)) /* synthesis syn_module_defined=1 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(32[13:44])
    inverter_U25 \inverter_chain_977..inv  (.\notGate[976]_keep (notGate_976), 
            .\notGate[977] (notGate_977)) /* synthesis syn_module_defined=1 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(32[13:44])
    inverter_U26 \inverter_chain_976..inv  (.\notGate[975]_keep (notGate_975), 
            .\notGate[976] (notGate_976)) /* synthesis syn_module_defined=1 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(32[13:44])
    inverter_U27 \inverter_chain_975..inv  (.\notGate[974]_keep (notGate_974), 
            .\notGate[975] (notGate_975)) /* synthesis syn_module_defined=1 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(32[13:44])
    inverter_U28 \inverter_chain_974..inv  (.\notGate[973]_keep (notGate_973), 
            .\notGate[974] (notGate_974)) /* synthesis syn_module_defined=1 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(32[13:44])
    inverter_U29 \inverter_chain_973..inv  (.\notGate[972]_keep (notGate_972), 
            .\notGate[973] (notGate_973)) /* synthesis syn_module_defined=1 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(32[13:44])
    inverter_U30 \inverter_chain_972..inv  (.\notGate[971]_keep (notGate_971), 
            .\notGate[972] (notGate_972)) /* synthesis syn_module_defined=1 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(32[13:44])
    inverter_U31 \inverter_chain_971..inv  (.\notGate[970]_keep (notGate_970), 
            .\notGate[971] (notGate_971)) /* synthesis syn_module_defined=1 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(32[13:44])
    inverter_U32 \inverter_chain_970..inv  (.\notGate[969]_keep (notGate_969), 
            .\notGate[970] (notGate_970)) /* synthesis syn_module_defined=1 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(32[13:44])
    inverter_U33 \inverter_chain_96..inv  (.\notGate[95]_keep (notGate_95), 
            .\notGate[96] (notGate_96)) /* synthesis syn_module_defined=1 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(32[13:44])
    inverter_U34 \inverter_chain_969..inv  (.\notGate[968]_keep (notGate_968), 
            .\notGate[969] (notGate_969)) /* synthesis syn_module_defined=1 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(32[13:44])
    inverter_U35 \inverter_chain_968..inv  (.\notGate[967]_keep (notGate_967), 
            .\notGate[968] (notGate_968)) /* synthesis syn_module_defined=1 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(32[13:44])
    inverter_U36 \inverter_chain_967..inv  (.\notGate[966]_keep (notGate_966), 
            .\notGate[967] (notGate_967)) /* synthesis syn_module_defined=1 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(32[13:44])
    inverter_U37 \inverter_chain_966..inv  (.\notGate[965]_keep (notGate_965), 
            .\notGate[966] (notGate_966)) /* synthesis syn_module_defined=1 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(32[13:44])
    inverter_U38 \inverter_chain_965..inv  (.\notGate[964]_keep (notGate_964), 
            .\notGate[965] (notGate_965)) /* synthesis syn_module_defined=1 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(32[13:44])
    inverter_U39 \inverter_chain_964..inv  (.\notGate[963]_keep (notGate_963), 
            .\notGate[964] (notGate_964)) /* synthesis syn_module_defined=1 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(32[13:44])
    inverter_U40 \inverter_chain_963..inv  (.\notGate[962]_keep (notGate_962), 
            .\notGate[963] (notGate_963)) /* synthesis syn_module_defined=1 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(32[13:44])
    inverter_U41 \inverter_chain_962..inv  (.\notGate[961]_keep (notGate_961), 
            .\notGate[962] (notGate_962)) /* synthesis syn_module_defined=1 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(32[13:44])
    inverter_U42 \inverter_chain_961..inv  (.\notGate[960]_keep (notGate_960), 
            .\notGate[961] (notGate_961)) /* synthesis syn_module_defined=1 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(32[13:44])
    inverter_U43 \inverter_chain_960..inv  (.\notGate[959]_keep (notGate_959), 
            .\notGate[960] (notGate_960)) /* synthesis syn_module_defined=1 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(32[13:44])
    inverter_U44 \inverter_chain_95..inv  (.\notGate[94]_keep (notGate_94), 
            .\notGate[95] (notGate_95)) /* synthesis syn_module_defined=1 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(32[13:44])
    inverter_U45 \inverter_chain_959..inv  (.\notGate[958]_keep (notGate_958), 
            .\notGate[959] (notGate_959)) /* synthesis syn_module_defined=1 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(32[13:44])
    inverter_U46 \inverter_chain_958..inv  (.\notGate[957]_keep (notGate_957), 
            .\notGate[958] (notGate_958)) /* synthesis syn_module_defined=1 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(32[13:44])
    inverter_U47 \inverter_chain_957..inv  (.\notGate[956]_keep (notGate_956), 
            .\notGate[957] (notGate_957)) /* synthesis syn_module_defined=1 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(32[13:44])
    inverter_U48 \inverter_chain_956..inv  (.\notGate[955]_keep (notGate_955), 
            .\notGate[956] (notGate_956)) /* synthesis syn_module_defined=1 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(32[13:44])
    inverter_U49 \inverter_chain_955..inv  (.\notGate[954]_keep (notGate_954), 
            .\notGate[955] (notGate_955)) /* synthesis syn_module_defined=1 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(32[13:44])
    inverter_U50 \inverter_chain_954..inv  (.\notGate[953]_keep (notGate_953), 
            .\notGate[954] (notGate_954)) /* synthesis syn_module_defined=1 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(32[13:44])
    inverter_U51 \inverter_chain_953..inv  (.\notGate[952]_keep (notGate_952), 
            .\notGate[953] (notGate_953)) /* synthesis syn_module_defined=1 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(32[13:44])
    inverter_U52 \inverter_chain_952..inv  (.\notGate[951]_keep (notGate_951), 
            .\notGate[952] (notGate_952)) /* synthesis syn_module_defined=1 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(32[13:44])
    inverter_U53 \inverter_chain_951..inv  (.\notGate[950]_keep (notGate_950), 
            .\notGate[951] (notGate_951)) /* synthesis syn_module_defined=1 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(32[13:44])
    inverter_U54 \inverter_chain_950..inv  (.\notGate[949]_keep (notGate_949), 
            .\notGate[950] (notGate_950)) /* synthesis syn_module_defined=1 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(32[13:44])
    inverter_U55 \inverter_chain_94..inv  (.\notGate[93]_keep (notGate_93), 
            .\notGate[94] (notGate_94)) /* synthesis syn_module_defined=1 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(32[13:44])
    inverter_U56 \inverter_chain_949..inv  (.\notGate[948]_keep (notGate_948), 
            .\notGate[949] (notGate_949)) /* synthesis syn_module_defined=1 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(32[13:44])
    inverter_U57 \inverter_chain_948..inv  (.\notGate[947]_keep (notGate_947), 
            .\notGate[948] (notGate_948)) /* synthesis syn_module_defined=1 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(32[13:44])
    inverter_U58 \inverter_chain_947..inv  (.\notGate[946]_keep (notGate_946), 
            .\notGate[947] (notGate_947)) /* synthesis syn_module_defined=1 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(32[13:44])
    inverter_U59 \inverter_chain_946..inv  (.\notGate[945]_keep (notGate_945), 
            .\notGate[946] (notGate_946)) /* synthesis syn_module_defined=1 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(32[13:44])
    inverter_U60 \inverter_chain_945..inv  (.\notGate[944]_keep (notGate_944), 
            .\notGate[945] (notGate_945)) /* synthesis syn_module_defined=1 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(32[13:44])
    inverter_U61 \inverter_chain_944..inv  (.\notGate[943]_keep (notGate_943), 
            .\notGate[944] (notGate_944)) /* synthesis syn_module_defined=1 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(32[13:44])
    inverter_U62 \inverter_chain_943..inv  (.\notGate[942]_keep (notGate_942), 
            .\notGate[943] (notGate_943)) /* synthesis syn_module_defined=1 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(32[13:44])
    inverter_U63 \inverter_chain_942..inv  (.\notGate[941]_keep (notGate_941), 
            .\notGate[942] (notGate_942)) /* synthesis syn_module_defined=1 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(32[13:44])
    inverter_U64 \inverter_chain_941..inv  (.\notGate[940]_keep (notGate_940), 
            .\notGate[941] (notGate_941)) /* synthesis syn_module_defined=1 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(32[13:44])
    inverter_U65 \inverter_chain_940..inv  (.\notGate[939]_keep (notGate_939), 
            .\notGate[940] (notGate_940)) /* synthesis syn_module_defined=1 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(32[13:44])
    inverter_U66 \inverter_chain_93..inv  (.\notGate[92]_keep (notGate_92), 
            .\notGate[93] (notGate_93)) /* synthesis syn_module_defined=1 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(32[13:44])
    inverter_U67 \inverter_chain_939..inv  (.\notGate[938]_keep (notGate_938), 
            .\notGate[939] (notGate_939)) /* synthesis syn_module_defined=1 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(32[13:44])
    inverter_U68 \inverter_chain_938..inv  (.\notGate[937]_keep (notGate_937), 
            .\notGate[938] (notGate_938)) /* synthesis syn_module_defined=1 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(32[13:44])
    inverter_U69 \inverter_chain_937..inv  (.\notGate[936]_keep (notGate_936), 
            .\notGate[937] (notGate_937)) /* synthesis syn_module_defined=1 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(32[13:44])
    inverter_U70 \inverter_chain_936..inv  (.\notGate[935]_keep (notGate_935), 
            .\notGate[936] (notGate_936)) /* synthesis syn_module_defined=1 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(32[13:44])
    inverter_U71 \inverter_chain_935..inv  (.\notGate[934]_keep (notGate_934), 
            .\notGate[935] (notGate_935)) /* synthesis syn_module_defined=1 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(32[13:44])
    inverter_U72 \inverter_chain_934..inv  (.\notGate[933]_keep (notGate_933), 
            .\notGate[934] (notGate_934)) /* synthesis syn_module_defined=1 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(32[13:44])
    inverter_U73 \inverter_chain_933..inv  (.\notGate[932]_keep (notGate_932), 
            .\notGate[933] (notGate_933)) /* synthesis syn_module_defined=1 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(32[13:44])
    inverter_U74 \inverter_chain_932..inv  (.\notGate[931]_keep (notGate_931), 
            .\notGate[932] (notGate_932)) /* synthesis syn_module_defined=1 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(32[13:44])
    inverter_U75 \inverter_chain_931..inv  (.\notGate[930]_keep (notGate_930), 
            .\notGate[931] (notGate_931)) /* synthesis syn_module_defined=1 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(32[13:44])
    inverter_U76 \inverter_chain_930..inv  (.\notGate[929]_keep (notGate_929), 
            .\notGate[930] (notGate_930)) /* synthesis syn_module_defined=1 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(32[13:44])
    inverter_U77 \inverter_chain_92..inv  (.\notGate[91]_keep (notGate_91), 
            .\notGate[92] (notGate_92)) /* synthesis syn_module_defined=1 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(32[13:44])
    inverter_U78 \inverter_chain_929..inv  (.\notGate[928]_keep (notGate_928), 
            .\notGate[929] (notGate_929)) /* synthesis syn_module_defined=1 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(32[13:44])
    inverter_U79 \inverter_chain_928..inv  (.\notGate[927]_keep (notGate_927), 
            .\notGate[928] (notGate_928)) /* synthesis syn_module_defined=1 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(32[13:44])
    inverter_U80 \inverter_chain_927..inv  (.\notGate[926]_keep (notGate_926), 
            .\notGate[927] (notGate_927)) /* synthesis syn_module_defined=1 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(32[13:44])
    inverter_U81 \inverter_chain_926..inv  (.\notGate[925]_keep (notGate_925), 
            .\notGate[926] (notGate_926)) /* synthesis syn_module_defined=1 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(32[13:44])
    inverter_U82 \inverter_chain_925..inv  (.\notGate[924]_keep (notGate_924), 
            .\notGate[925] (notGate_925)) /* synthesis syn_module_defined=1 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(32[13:44])
    inverter_U83 \inverter_chain_924..inv  (.\notGate[923]_keep (notGate_923), 
            .\notGate[924] (notGate_924)) /* synthesis syn_module_defined=1 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(32[13:44])
    inverter_U84 \inverter_chain_923..inv  (.\notGate[922]_keep (notGate_922), 
            .\notGate[923] (notGate_923)) /* synthesis syn_module_defined=1 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(32[13:44])
    inverter_U85 \inverter_chain_922..inv  (.\notGate[921]_keep (notGate_921), 
            .\notGate[922] (notGate_922)) /* synthesis syn_module_defined=1 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(32[13:44])
    inverter_U86 \inverter_chain_921..inv  (.\notGate[920]_keep (notGate_920), 
            .\notGate[921] (notGate_921)) /* synthesis syn_module_defined=1 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(32[13:44])
    inverter_U87 \inverter_chain_920..inv  (.\notGate[919]_keep (notGate_919), 
            .\notGate[920] (notGate_920)) /* synthesis syn_module_defined=1 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(32[13:44])
    inverter_U88 \inverter_chain_91..inv  (.\notGate[90]_keep (notGate_90), 
            .\notGate[91] (notGate_91)) /* synthesis syn_module_defined=1 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(32[13:44])
    inverter_U89 \inverter_chain_919..inv  (.\notGate[918]_keep (notGate_918), 
            .\notGate[919] (notGate_919)) /* synthesis syn_module_defined=1 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(32[13:44])
    inverter_U90 \inverter_chain_918..inv  (.\notGate[917]_keep (notGate_917), 
            .\notGate[918] (notGate_918)) /* synthesis syn_module_defined=1 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(32[13:44])
    inverter_U91 \inverter_chain_917..inv  (.\notGate[916]_keep (notGate_916), 
            .\notGate[917] (notGate_917)) /* synthesis syn_module_defined=1 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(32[13:44])
    inverter_U92 \inverter_chain_916..inv  (.\notGate[915]_keep (notGate_915), 
            .\notGate[916] (notGate_916)) /* synthesis syn_module_defined=1 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(32[13:44])
    inverter_U93 \inverter_chain_915..inv  (.\notGate[914]_keep (notGate_914), 
            .\notGate[915] (notGate_915)) /* synthesis syn_module_defined=1 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(32[13:44])
    inverter_U94 \inverter_chain_914..inv  (.\notGate[913]_keep (notGate_913), 
            .\notGate[914] (notGate_914)) /* synthesis syn_module_defined=1 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(32[13:44])
    inverter_U95 \inverter_chain_913..inv  (.\notGate[912]_keep (notGate_912), 
            .\notGate[913] (notGate_913)) /* synthesis syn_module_defined=1 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(32[13:44])
    inverter_U96 \inverter_chain_912..inv  (.\notGate[911]_keep (notGate_911), 
            .\notGate[912] (notGate_912)) /* synthesis syn_module_defined=1 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(32[13:44])
    inverter_U97 \inverter_chain_911..inv  (.\notGate[910]_keep (notGate_910), 
            .\notGate[911] (notGate_911)) /* synthesis syn_module_defined=1 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(32[13:44])
    inverter_U98 \inverter_chain_910..inv  (.\notGate[909]_keep (notGate_909), 
            .\notGate[910] (notGate_910)) /* synthesis syn_module_defined=1 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(32[13:44])
    inverter_U99 \inverter_chain_90..inv  (.\notGate[89]_keep (notGate_89), 
            .\notGate[90] (notGate_90)) /* synthesis syn_module_defined=1 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(32[13:44])
    inverter_U100 \inverter_chain_909..inv  (.\notGate[908]_keep (notGate_908), 
            .\notGate[909] (notGate_909)) /* synthesis syn_module_defined=1 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(32[13:44])
    inverter_U101 \inverter_chain_908..inv  (.\notGate[907]_keep (notGate_907), 
            .\notGate[908] (notGate_908)) /* synthesis syn_module_defined=1 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(32[13:44])
    inverter_U102 \inverter_chain_907..inv  (.\notGate[906]_keep (notGate_906), 
            .\notGate[907] (notGate_907)) /* synthesis syn_module_defined=1 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(32[13:44])
    inverter_U103 \inverter_chain_906..inv  (.\notGate[905]_keep (notGate_905), 
            .\notGate[906] (notGate_906)) /* synthesis syn_module_defined=1 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(32[13:44])
    inverter_U104 \inverter_chain_905..inv  (.\notGate[904]_keep (notGate_904), 
            .\notGate[905] (notGate_905)) /* synthesis syn_module_defined=1 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(32[13:44])
    inverter_U105 \inverter_chain_904..inv  (.\notGate[903]_keep (notGate_903), 
            .\notGate[904] (notGate_904)) /* synthesis syn_module_defined=1 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(32[13:44])
    inverter_U106 \inverter_chain_903..inv  (.\notGate[902]_keep (notGate_902), 
            .\notGate[903] (notGate_903)) /* synthesis syn_module_defined=1 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(32[13:44])
    inverter_U107 \inverter_chain_902..inv  (.\notGate[901]_keep (notGate_901), 
            .\notGate[902] (notGate_902)) /* synthesis syn_module_defined=1 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(32[13:44])
    inverter_U108 \inverter_chain_901..inv  (.\notGate[900]_keep (notGate_900), 
            .\notGate[901] (notGate_901)) /* synthesis syn_module_defined=1 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(32[13:44])
    inverter_U109 \inverter_chain_900..inv  (.\notGate[899]_keep (notGate_899), 
            .\notGate[900] (notGate_900)) /* synthesis syn_module_defined=1 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(32[13:44])
    inverter_U110 \inverter_chain_8..inv  (.\notGate[7]_keep (notGate_7), 
            .\notGate[8] (notGate_8)) /* synthesis syn_module_defined=1 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(32[13:44])
    inverter_U111 \inverter_chain_89..inv  (.\notGate[88]_keep (notGate_88), 
            .\notGate[89] (notGate_89)) /* synthesis syn_module_defined=1 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(32[13:44])
    inverter_U112 \inverter_chain_899..inv  (.\notGate[898]_keep (notGate_898), 
            .\notGate[899] (notGate_899)) /* synthesis syn_module_defined=1 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(32[13:44])
    inverter_U113 \inverter_chain_898..inv  (.\notGate[897]_keep (notGate_897), 
            .\notGate[898] (notGate_898)) /* synthesis syn_module_defined=1 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(32[13:44])
    inverter_U114 \inverter_chain_897..inv  (.\notGate[896]_keep (notGate_896), 
            .\notGate[897] (notGate_897)) /* synthesis syn_module_defined=1 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(32[13:44])
    inverter_U115 \inverter_chain_896..inv  (.\notGate[895]_keep (notGate_895), 
            .\notGate[896] (notGate_896)) /* synthesis syn_module_defined=1 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(32[13:44])
    inverter_U116 \inverter_chain_895..inv  (.\notGate[894]_keep (notGate_894), 
            .\notGate[895] (notGate_895)) /* synthesis syn_module_defined=1 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(32[13:44])
    inverter_U117 \inverter_chain_894..inv  (.\notGate[893]_keep (notGate_893), 
            .\notGate[894] (notGate_894)) /* synthesis syn_module_defined=1 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(32[13:44])
    inverter_U118 \inverter_chain_893..inv  (.\notGate[892]_keep (notGate_892), 
            .\notGate[893] (notGate_893)) /* synthesis syn_module_defined=1 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(32[13:44])
    inverter_U119 \inverter_chain_892..inv  (.\notGate[891]_keep (notGate_891), 
            .\notGate[892] (notGate_892)) /* synthesis syn_module_defined=1 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(32[13:44])
    inverter_U120 \inverter_chain_891..inv  (.\notGate[890]_keep (notGate_890), 
            .\notGate[891] (notGate_891)) /* synthesis syn_module_defined=1 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(32[13:44])
    inverter_U121 \inverter_chain_890..inv  (.\notGate[889]_keep (notGate_889), 
            .\notGate[890] (notGate_890)) /* synthesis syn_module_defined=1 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(32[13:44])
    inverter_U122 \inverter_chain_88..inv  (.\notGate[87]_keep (notGate_87), 
            .\notGate[88] (notGate_88)) /* synthesis syn_module_defined=1 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(32[13:44])
    inverter_U123 \inverter_chain_889..inv  (.\notGate[888]_keep (notGate_888), 
            .\notGate[889] (notGate_889)) /* synthesis syn_module_defined=1 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(32[13:44])
    inverter_U124 \inverter_chain_888..inv  (.\notGate[887]_keep (notGate_887), 
            .\notGate[888] (notGate_888)) /* synthesis syn_module_defined=1 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(32[13:44])
    inverter_U125 \inverter_chain_887..inv  (.\notGate[886]_keep (notGate_886), 
            .\notGate[887] (notGate_887)) /* synthesis syn_module_defined=1 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(32[13:44])
    inverter_U126 \inverter_chain_886..inv  (.\notGate[885]_keep (notGate_885), 
            .\notGate[886] (notGate_886)) /* synthesis syn_module_defined=1 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(32[13:44])
    inverter_U127 \inverter_chain_885..inv  (.\notGate[884]_keep (notGate_884), 
            .\notGate[885] (notGate_885)) /* synthesis syn_module_defined=1 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(32[13:44])
    inverter_U128 \inverter_chain_884..inv  (.\notGate[883]_keep (notGate_883), 
            .\notGate[884] (notGate_884)) /* synthesis syn_module_defined=1 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(32[13:44])
    inverter_U129 \inverter_chain_883..inv  (.\notGate[882]_keep (notGate_882), 
            .\notGate[883] (notGate_883)) /* synthesis syn_module_defined=1 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(32[13:44])
    inverter_U130 \inverter_chain_882..inv  (.\notGate[881]_keep (notGate_881), 
            .\notGate[882] (notGate_882)) /* synthesis syn_module_defined=1 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(32[13:44])
    inverter_U131 \inverter_chain_881..inv  (.\notGate[880]_keep (notGate_880), 
            .\notGate[881] (notGate_881)) /* synthesis syn_module_defined=1 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(32[13:44])
    inverter_U132 \inverter_chain_880..inv  (.\notGate[879]_keep (notGate_879), 
            .\notGate[880] (notGate_880)) /* synthesis syn_module_defined=1 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(32[13:44])
    inverter_U133 \inverter_chain_87..inv  (.\notGate[86]_keep (notGate_86), 
            .\notGate[87] (notGate_87)) /* synthesis syn_module_defined=1 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(32[13:44])
    inverter_U134 \inverter_chain_879..inv  (.\notGate[878]_keep (notGate_878), 
            .\notGate[879] (notGate_879)) /* synthesis syn_module_defined=1 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(32[13:44])
    inverter_U135 \inverter_chain_878..inv  (.\notGate[877]_keep (notGate_877), 
            .\notGate[878] (notGate_878)) /* synthesis syn_module_defined=1 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(32[13:44])
    inverter_U136 \inverter_chain_877..inv  (.\notGate[876]_keep (notGate_876), 
            .\notGate[877] (notGate_877)) /* synthesis syn_module_defined=1 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(32[13:44])
    inverter_U137 \inverter_chain_876..inv  (.\notGate[875]_keep (notGate_875), 
            .\notGate[876] (notGate_876)) /* synthesis syn_module_defined=1 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(32[13:44])
    inverter_U138 \inverter_chain_875..inv  (.\notGate[874]_keep (notGate_874), 
            .\notGate[875] (notGate_875)) /* synthesis syn_module_defined=1 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(32[13:44])
    inverter_U139 \inverter_chain_874..inv  (.\notGate[873]_keep (notGate_873), 
            .\notGate[874] (notGate_874)) /* synthesis syn_module_defined=1 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(32[13:44])
    inverter_U140 \inverter_chain_873..inv  (.\notGate[872]_keep (notGate_872), 
            .\notGate[873] (notGate_873)) /* synthesis syn_module_defined=1 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(32[13:44])
    inverter_U141 \inverter_chain_872..inv  (.\notGate[871]_keep (notGate_871), 
            .\notGate[872] (notGate_872)) /* synthesis syn_module_defined=1 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(32[13:44])
    inverter_U142 \inverter_chain_871..inv  (.\notGate[870]_keep (notGate_870), 
            .\notGate[871] (notGate_871)) /* synthesis syn_module_defined=1 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(32[13:44])
    inverter_U143 \inverter_chain_870..inv  (.\notGate[869]_keep (notGate_869), 
            .\notGate[870] (notGate_870)) /* synthesis syn_module_defined=1 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(32[13:44])
    inverter_U144 \inverter_chain_86..inv  (.\notGate[85]_keep (notGate_85), 
            .\notGate[86] (notGate_86)) /* synthesis syn_module_defined=1 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(32[13:44])
    inverter_U145 \inverter_chain_869..inv  (.\notGate[868]_keep (notGate_868), 
            .\notGate[869] (notGate_869)) /* synthesis syn_module_defined=1 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(32[13:44])
    inverter_U146 \inverter_chain_868..inv  (.\notGate[867]_keep (notGate_867), 
            .\notGate[868] (notGate_868)) /* synthesis syn_module_defined=1 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(32[13:44])
    inverter_U147 \inverter_chain_867..inv  (.\notGate[866]_keep (notGate_866), 
            .\notGate[867] (notGate_867)) /* synthesis syn_module_defined=1 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(32[13:44])
    inverter_U148 \inverter_chain_866..inv  (.\notGate[865]_keep (notGate_865), 
            .\notGate[866] (notGate_866)) /* synthesis syn_module_defined=1 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(32[13:44])
    inverter_U149 \inverter_chain_865..inv  (.\notGate[864]_keep (notGate_864), 
            .\notGate[865] (notGate_865)) /* synthesis syn_module_defined=1 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(32[13:44])
    inverter_U150 \inverter_chain_864..inv  (.\notGate[863]_keep (notGate_863), 
            .\notGate[864] (notGate_864)) /* synthesis syn_module_defined=1 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(32[13:44])
    inverter_U151 \inverter_chain_863..inv  (.\notGate[862]_keep (notGate_862), 
            .\notGate[863] (notGate_863)) /* synthesis syn_module_defined=1 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(32[13:44])
    inverter_U152 \inverter_chain_862..inv  (.\notGate[861]_keep (notGate_861), 
            .\notGate[862] (notGate_862)) /* synthesis syn_module_defined=1 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(32[13:44])
    inverter_U153 \inverter_chain_861..inv  (.\notGate[860]_keep (notGate_860), 
            .\notGate[861] (notGate_861)) /* synthesis syn_module_defined=1 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(32[13:44])
    inverter_U154 \inverter_chain_860..inv  (.\notGate[859]_keep (notGate_859), 
            .\notGate[860] (notGate_860)) /* synthesis syn_module_defined=1 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(32[13:44])
    inverter_U155 \inverter_chain_85..inv  (.\notGate[84]_keep (notGate_84), 
            .\notGate[85] (notGate_85)) /* synthesis syn_module_defined=1 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(32[13:44])
    inverter_U156 \inverter_chain_859..inv  (.\notGate[858]_keep (notGate_858), 
            .\notGate[859] (notGate_859)) /* synthesis syn_module_defined=1 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(32[13:44])
    inverter_U157 \inverter_chain_858..inv  (.\notGate[857]_keep (notGate_857), 
            .\notGate[858] (notGate_858)) /* synthesis syn_module_defined=1 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(32[13:44])
    inverter_U158 \inverter_chain_857..inv  (.\notGate[856]_keep (notGate_856), 
            .\notGate[857] (notGate_857)) /* synthesis syn_module_defined=1 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(32[13:44])
    inverter_U159 \inverter_chain_856..inv  (.\notGate[855]_keep (notGate_855), 
            .\notGate[856] (notGate_856)) /* synthesis syn_module_defined=1 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(32[13:44])
    inverter_U160 \inverter_chain_855..inv  (.\notGate[854]_keep (notGate_854), 
            .\notGate[855] (notGate_855)) /* synthesis syn_module_defined=1 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(32[13:44])
    inverter_U161 \inverter_chain_854..inv  (.\notGate[853]_keep (notGate_853), 
            .\notGate[854] (notGate_854)) /* synthesis syn_module_defined=1 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(32[13:44])
    inverter_U162 \inverter_chain_853..inv  (.\notGate[852]_keep (notGate_852), 
            .\notGate[853] (notGate_853)) /* synthesis syn_module_defined=1 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(32[13:44])
    inverter_U163 \inverter_chain_852..inv  (.\notGate[851]_keep (notGate_851), 
            .\notGate[852] (notGate_852)) /* synthesis syn_module_defined=1 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(32[13:44])
    inverter_U164 \inverter_chain_851..inv  (.\notGate[850]_keep (notGate_850), 
            .\notGate[851] (notGate_851)) /* synthesis syn_module_defined=1 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(32[13:44])
    inverter_U165 \inverter_chain_850..inv  (.\notGate[849]_keep (notGate_849), 
            .\notGate[850] (notGate_850)) /* synthesis syn_module_defined=1 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(32[13:44])
    inverter_U166 \inverter_chain_84..inv  (.\notGate[83]_keep (notGate_83), 
            .\notGate[84] (notGate_84)) /* synthesis syn_module_defined=1 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(32[13:44])
    inverter_U167 \inverter_chain_849..inv  (.\notGate[848]_keep (notGate_848), 
            .\notGate[849] (notGate_849)) /* synthesis syn_module_defined=1 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(32[13:44])
    inverter_U168 \inverter_chain_848..inv  (.\notGate[847]_keep (notGate_847), 
            .\notGate[848] (notGate_848)) /* synthesis syn_module_defined=1 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(32[13:44])
    inverter_U169 \inverter_chain_847..inv  (.\notGate[846]_keep (notGate_846), 
            .\notGate[847] (notGate_847)) /* synthesis syn_module_defined=1 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(32[13:44])
    inverter_U170 \inverter_chain_846..inv  (.\notGate[845]_keep (notGate_845), 
            .\notGate[846] (notGate_846)) /* synthesis syn_module_defined=1 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(32[13:44])
    inverter_U171 \inverter_chain_845..inv  (.\notGate[844]_keep (notGate_844), 
            .\notGate[845] (notGate_845)) /* synthesis syn_module_defined=1 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(32[13:44])
    inverter_U172 \inverter_chain_844..inv  (.\notGate[843]_keep (notGate_843), 
            .\notGate[844] (notGate_844)) /* synthesis syn_module_defined=1 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(32[13:44])
    inverter_U173 \inverter_chain_843..inv  (.\notGate[842]_keep (notGate_842), 
            .\notGate[843] (notGate_843)) /* synthesis syn_module_defined=1 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(32[13:44])
    inverter_U174 \inverter_chain_842..inv  (.\notGate[841]_keep (notGate_841), 
            .\notGate[842] (notGate_842)) /* synthesis syn_module_defined=1 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(32[13:44])
    inverter_U175 \inverter_chain_841..inv  (.\notGate[840]_keep (notGate_840), 
            .\notGate[841] (notGate_841)) /* synthesis syn_module_defined=1 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(32[13:44])
    inverter_U176 \inverter_chain_840..inv  (.\notGate[839]_keep (notGate_839), 
            .\notGate[840] (notGate_840)) /* synthesis syn_module_defined=1 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(32[13:44])
    inverter_U177 \inverter_chain_83..inv  (.\notGate[82]_keep (notGate_82), 
            .\notGate[83] (notGate_83)) /* synthesis syn_module_defined=1 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(32[13:44])
    inverter_U178 \inverter_chain_839..inv  (.\notGate[838]_keep (notGate_838), 
            .\notGate[839] (notGate_839)) /* synthesis syn_module_defined=1 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(32[13:44])
    inverter_U179 \inverter_chain_838..inv  (.\notGate[837]_keep (notGate_837), 
            .\notGate[838] (notGate_838)) /* synthesis syn_module_defined=1 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(32[13:44])
    inverter_U180 \inverter_chain_837..inv  (.\notGate[836]_keep (notGate_836), 
            .\notGate[837] (notGate_837)) /* synthesis syn_module_defined=1 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(32[13:44])
    inverter_U181 \inverter_chain_836..inv  (.\notGate[835]_keep (notGate_835), 
            .\notGate[836] (notGate_836)) /* synthesis syn_module_defined=1 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(32[13:44])
    inverter_U182 \inverter_chain_835..inv  (.\notGate[834]_keep (notGate_834), 
            .\notGate[835] (notGate_835)) /* synthesis syn_module_defined=1 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(32[13:44])
    inverter_U183 \inverter_chain_834..inv  (.\notGate[833]_keep (notGate_833), 
            .\notGate[834] (notGate_834)) /* synthesis syn_module_defined=1 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(32[13:44])
    inverter_U184 \inverter_chain_833..inv  (.\notGate[832]_keep (notGate_832), 
            .\notGate[833] (notGate_833)) /* synthesis syn_module_defined=1 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(32[13:44])
    inverter_U185 \inverter_chain_832..inv  (.\notGate[831]_keep (notGate_831), 
            .\notGate[832] (notGate_832)) /* synthesis syn_module_defined=1 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(32[13:44])
    inverter_U186 \inverter_chain_831..inv  (.\notGate[830]_keep (notGate_830), 
            .\notGate[831] (notGate_831)) /* synthesis syn_module_defined=1 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(32[13:44])
    inverter_U187 \inverter_chain_830..inv  (.\notGate[829]_keep (notGate_829), 
            .\notGate[830] (notGate_830)) /* synthesis syn_module_defined=1 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(32[13:44])
    inverter_U188 \inverter_chain_82..inv  (.\notGate[81]_keep (notGate_81), 
            .\notGate[82] (notGate_82)) /* synthesis syn_module_defined=1 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(32[13:44])
    inverter_U189 \inverter_chain_829..inv  (.\notGate[828]_keep (notGate_828), 
            .\notGate[829] (notGate_829)) /* synthesis syn_module_defined=1 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(32[13:44])
    inverter_U190 \inverter_chain_828..inv  (.\notGate[827]_keep (notGate_827), 
            .\notGate[828] (notGate_828)) /* synthesis syn_module_defined=1 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(32[13:44])
    inverter_U191 \inverter_chain_827..inv  (.\notGate[826]_keep (notGate_826), 
            .\notGate[827] (notGate_827)) /* synthesis syn_module_defined=1 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(32[13:44])
    inverter_U192 \inverter_chain_826..inv  (.\notGate[825]_keep (notGate_825), 
            .\notGate[826] (notGate_826)) /* synthesis syn_module_defined=1 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(32[13:44])
    inverter_U193 \inverter_chain_825..inv  (.\notGate[824]_keep (notGate_824), 
            .\notGate[825] (notGate_825)) /* synthesis syn_module_defined=1 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(32[13:44])
    inverter_U194 \inverter_chain_824..inv  (.\notGate[823]_keep (notGate_823), 
            .\notGate[824] (notGate_824)) /* synthesis syn_module_defined=1 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(32[13:44])
    inverter_U195 \inverter_chain_823..inv  (.\notGate[822]_keep (notGate_822), 
            .\notGate[823] (notGate_823)) /* synthesis syn_module_defined=1 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(32[13:44])
    inverter_U196 \inverter_chain_822..inv  (.\notGate[821]_keep (notGate_821), 
            .\notGate[822] (notGate_822)) /* synthesis syn_module_defined=1 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(32[13:44])
    inverter_U197 \inverter_chain_821..inv  (.\notGate[820]_keep (notGate_820), 
            .\notGate[821] (notGate_821)) /* synthesis syn_module_defined=1 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(32[13:44])
    inverter_U198 \inverter_chain_820..inv  (.\notGate[819]_keep (notGate_819), 
            .\notGate[820] (notGate_820)) /* synthesis syn_module_defined=1 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(32[13:44])
    inverter_U199 \inverter_chain_81..inv  (.\notGate[80]_keep (notGate_80), 
            .\notGate[81] (notGate_81)) /* synthesis syn_module_defined=1 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(32[13:44])
    inverter_U200 \inverter_chain_819..inv  (.\notGate[818]_keep (notGate_818), 
            .\notGate[819] (notGate_819)) /* synthesis syn_module_defined=1 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(32[13:44])
    inverter_U201 \inverter_chain_818..inv  (.\notGate[817]_keep (notGate_817), 
            .\notGate[818] (notGate_818)) /* synthesis syn_module_defined=1 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(32[13:44])
    inverter_U202 \inverter_chain_817..inv  (.\notGate[816]_keep (notGate_816), 
            .\notGate[817] (notGate_817)) /* synthesis syn_module_defined=1 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(32[13:44])
    inverter_U203 \inverter_chain_816..inv  (.\notGate[815]_keep (notGate_815), 
            .\notGate[816] (notGate_816)) /* synthesis syn_module_defined=1 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(32[13:44])
    inverter_U204 \inverter_chain_815..inv  (.\notGate[814]_keep (notGate_814), 
            .\notGate[815] (notGate_815)) /* synthesis syn_module_defined=1 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(32[13:44])
    inverter_U205 \inverter_chain_814..inv  (.\notGate[813]_keep (notGate_813), 
            .\notGate[814] (notGate_814)) /* synthesis syn_module_defined=1 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(32[13:44])
    inverter_U206 \inverter_chain_813..inv  (.\notGate[812]_keep (notGate_812), 
            .\notGate[813] (notGate_813)) /* synthesis syn_module_defined=1 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(32[13:44])
    inverter_U207 \inverter_chain_812..inv  (.\notGate[811]_keep (notGate_811), 
            .\notGate[812] (notGate_812)) /* synthesis syn_module_defined=1 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(32[13:44])
    inverter_U208 \inverter_chain_811..inv  (.\notGate[810]_keep (notGate_810), 
            .\notGate[811] (notGate_811)) /* synthesis syn_module_defined=1 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(32[13:44])
    inverter_U209 \inverter_chain_810..inv  (.\notGate[809]_keep (notGate_809), 
            .\notGate[810] (notGate_810)) /* synthesis syn_module_defined=1 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(32[13:44])
    inverter_U210 \inverter_chain_80..inv  (.\notGate[79]_keep (notGate_79), 
            .\notGate[80] (notGate_80)) /* synthesis syn_module_defined=1 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(32[13:44])
    inverter_U211 \inverter_chain_809..inv  (.\notGate[808]_keep (notGate_808), 
            .\notGate[809] (notGate_809)) /* synthesis syn_module_defined=1 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(32[13:44])
    inverter_U212 \inverter_chain_808..inv  (.\notGate[807]_keep (notGate_807), 
            .\notGate[808] (notGate_808)) /* synthesis syn_module_defined=1 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(32[13:44])
    inverter_U213 \inverter_chain_807..inv  (.\notGate[806]_keep (notGate_806), 
            .\notGate[807] (notGate_807)) /* synthesis syn_module_defined=1 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(32[13:44])
    inverter_U214 \inverter_chain_806..inv  (.\notGate[805]_keep (notGate_805), 
            .\notGate[806] (notGate_806)) /* synthesis syn_module_defined=1 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(32[13:44])
    inverter_U215 \inverter_chain_805..inv  (.\notGate[804]_keep (notGate_804), 
            .\notGate[805] (notGate_805)) /* synthesis syn_module_defined=1 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(32[13:44])
    inverter_U216 \inverter_chain_804..inv  (.\notGate[803]_keep (notGate_803), 
            .\notGate[804] (notGate_804)) /* synthesis syn_module_defined=1 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(32[13:44])
    inverter_U217 \inverter_chain_803..inv  (.\notGate[802]_keep (notGate_802), 
            .\notGate[803] (notGate_803)) /* synthesis syn_module_defined=1 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(32[13:44])
    inverter_U218 \inverter_chain_802..inv  (.\notGate[801]_keep (notGate_801), 
            .\notGate[802] (notGate_802)) /* synthesis syn_module_defined=1 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(32[13:44])
    inverter_U219 \inverter_chain_801..inv  (.\notGate[800]_keep (notGate_800), 
            .\notGate[801] (notGate_801)) /* synthesis syn_module_defined=1 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(32[13:44])
    inverter_U220 \inverter_chain_800..inv  (.\notGate[799]_keep (notGate_799), 
            .\notGate[800] (notGate_800)) /* synthesis syn_module_defined=1 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(32[13:44])
    inverter_U221 \inverter_chain_7..inv  (.\notGate[6]_keep (notGate_6), 
            .\notGate[7] (notGate_7)) /* synthesis syn_module_defined=1 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(32[13:44])
    inverter_U222 \inverter_chain_79..inv  (.\notGate[78]_keep (notGate_78), 
            .\notGate[79] (notGate_79)) /* synthesis syn_module_defined=1 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(32[13:44])
    inverter_U223 \inverter_chain_799..inv  (.\notGate[798]_keep (notGate_798), 
            .\notGate[799] (notGate_799)) /* synthesis syn_module_defined=1 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(32[13:44])
    inverter_U224 \inverter_chain_798..inv  (.\notGate[797]_keep (notGate_797), 
            .\notGate[798] (notGate_798)) /* synthesis syn_module_defined=1 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(32[13:44])
    inverter_U225 \inverter_chain_797..inv  (.\notGate[796]_keep (notGate_796), 
            .\notGate[797] (notGate_797)) /* synthesis syn_module_defined=1 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(32[13:44])
    inverter_U226 \inverter_chain_796..inv  (.\notGate[795]_keep (notGate_795), 
            .\notGate[796] (notGate_796)) /* synthesis syn_module_defined=1 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(32[13:44])
    inverter_U227 \inverter_chain_795..inv  (.\notGate[794]_keep (notGate_794), 
            .\notGate[795] (notGate_795)) /* synthesis syn_module_defined=1 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(32[13:44])
    inverter_U228 \inverter_chain_794..inv  (.\notGate[793]_keep (notGate_793), 
            .\notGate[794] (notGate_794)) /* synthesis syn_module_defined=1 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(32[13:44])
    inverter_U229 \inverter_chain_793..inv  (.\notGate[792]_keep (notGate_792), 
            .\notGate[793] (notGate_793)) /* synthesis syn_module_defined=1 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(32[13:44])
    inverter_U230 \inverter_chain_792..inv  (.\notGate[791]_keep (notGate_791), 
            .\notGate[792] (notGate_792)) /* synthesis syn_module_defined=1 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(32[13:44])
    inverter_U231 \inverter_chain_791..inv  (.\notGate[790]_keep (notGate_790), 
            .\notGate[791] (notGate_791)) /* synthesis syn_module_defined=1 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(32[13:44])
    inverter_U232 \inverter_chain_790..inv  (.\notGate[789]_keep (notGate_789), 
            .\notGate[790] (notGate_790)) /* synthesis syn_module_defined=1 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(32[13:44])
    inverter_U233 \inverter_chain_78..inv  (.\notGate[77]_keep (notGate_77), 
            .\notGate[78] (notGate_78)) /* synthesis syn_module_defined=1 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(32[13:44])
    inverter_U234 \inverter_chain_789..inv  (.\notGate[788]_keep (notGate_788), 
            .\notGate[789] (notGate_789)) /* synthesis syn_module_defined=1 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(32[13:44])
    inverter_U235 \inverter_chain_788..inv  (.\notGate[787]_keep (notGate_787), 
            .\notGate[788] (notGate_788)) /* synthesis syn_module_defined=1 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(32[13:44])
    inverter_U236 \inverter_chain_787..inv  (.\notGate[786]_keep (notGate_786), 
            .\notGate[787] (notGate_787)) /* synthesis syn_module_defined=1 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(32[13:44])
    inverter_U237 \inverter_chain_786..inv  (.\notGate[785]_keep (notGate_785), 
            .\notGate[786] (notGate_786)) /* synthesis syn_module_defined=1 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(32[13:44])
    inverter_U238 \inverter_chain_785..inv  (.\notGate[784]_keep (notGate_784), 
            .\notGate[785] (notGate_785)) /* synthesis syn_module_defined=1 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(32[13:44])
    inverter_U239 \inverter_chain_784..inv  (.\notGate[783]_keep (notGate_783), 
            .\notGate[784] (notGate_784)) /* synthesis syn_module_defined=1 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(32[13:44])
    inverter_U240 \inverter_chain_783..inv  (.\notGate[782]_keep (notGate_782), 
            .\notGate[783] (notGate_783)) /* synthesis syn_module_defined=1 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(32[13:44])
    inverter_U241 \inverter_chain_782..inv  (.\notGate[781]_keep (notGate_781), 
            .\notGate[782] (notGate_782)) /* synthesis syn_module_defined=1 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(32[13:44])
    inverter_U242 \inverter_chain_781..inv  (.\notGate[780]_keep (notGate_780), 
            .\notGate[781] (notGate_781)) /* synthesis syn_module_defined=1 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(32[13:44])
    inverter_U243 \inverter_chain_780..inv  (.\notGate[779]_keep (notGate_779), 
            .\notGate[780] (notGate_780)) /* synthesis syn_module_defined=1 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(32[13:44])
    inverter_U244 \inverter_chain_77..inv  (.\notGate[76]_keep (notGate_76), 
            .\notGate[77] (notGate_77)) /* synthesis syn_module_defined=1 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(32[13:44])
    inverter_U245 \inverter_chain_779..inv  (.\notGate[778]_keep (notGate_778), 
            .\notGate[779] (notGate_779)) /* synthesis syn_module_defined=1 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(32[13:44])
    inverter_U246 \inverter_chain_778..inv  (.\notGate[777]_keep (notGate_777), 
            .\notGate[778] (notGate_778)) /* synthesis syn_module_defined=1 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(32[13:44])
    inverter_U247 \inverter_chain_777..inv  (.\notGate[776]_keep (notGate_776), 
            .\notGate[777] (notGate_777)) /* synthesis syn_module_defined=1 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(32[13:44])
    inverter_U248 \inverter_chain_776..inv  (.\notGate[775]_keep (notGate_775), 
            .\notGate[776] (notGate_776)) /* synthesis syn_module_defined=1 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(32[13:44])
    inverter_U249 \inverter_chain_775..inv  (.\notGate[774]_keep (notGate_774), 
            .\notGate[775] (notGate_775)) /* synthesis syn_module_defined=1 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(32[13:44])
    inverter_U250 \inverter_chain_774..inv  (.\notGate[773]_keep (notGate_773), 
            .\notGate[774] (notGate_774)) /* synthesis syn_module_defined=1 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(32[13:44])
    inverter_U251 \inverter_chain_773..inv  (.\notGate[772]_keep (notGate_772), 
            .\notGate[773] (notGate_773)) /* synthesis syn_module_defined=1 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(32[13:44])
    inverter_U252 \inverter_chain_772..inv  (.\notGate[771]_keep (notGate_771), 
            .\notGate[772] (notGate_772)) /* synthesis syn_module_defined=1 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(32[13:44])
    inverter_U253 \inverter_chain_771..inv  (.\notGate[770]_keep (notGate_770), 
            .\notGate[771] (notGate_771)) /* synthesis syn_module_defined=1 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(32[13:44])
    inverter_U254 \inverter_chain_770..inv  (.\notGate[769]_keep (notGate_769), 
            .\notGate[770] (notGate_770)) /* synthesis syn_module_defined=1 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(32[13:44])
    inverter_U255 \inverter_chain_76..inv  (.\notGate[75]_keep (notGate_75), 
            .\notGate[76] (notGate_76)) /* synthesis syn_module_defined=1 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(32[13:44])
    inverter_U256 \inverter_chain_769..inv  (.\notGate[768]_keep (notGate_768), 
            .\notGate[769] (notGate_769)) /* synthesis syn_module_defined=1 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(32[13:44])
    inverter_U257 \inverter_chain_768..inv  (.\notGate[767]_keep (notGate_767), 
            .\notGate[768] (notGate_768)) /* synthesis syn_module_defined=1 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(32[13:44])
    inverter_U258 \inverter_chain_767..inv  (.\notGate[766]_keep (notGate_766), 
            .\notGate[767] (notGate_767)) /* synthesis syn_module_defined=1 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(32[13:44])
    inverter_U259 \inverter_chain_766..inv  (.\notGate[765]_keep (notGate_765), 
            .\notGate[766] (notGate_766)) /* synthesis syn_module_defined=1 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(32[13:44])
    inverter_U260 \inverter_chain_765..inv  (.\notGate[764]_keep (notGate_764), 
            .\notGate[765] (notGate_765)) /* synthesis syn_module_defined=1 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(32[13:44])
    inverter_U261 \inverter_chain_764..inv  (.\notGate[763]_keep (notGate_763), 
            .\notGate[764] (notGate_764)) /* synthesis syn_module_defined=1 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(32[13:44])
    inverter_U262 \inverter_chain_763..inv  (.\notGate[762]_keep (notGate_762), 
            .\notGate[763] (notGate_763)) /* synthesis syn_module_defined=1 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(32[13:44])
    inverter_U263 \inverter_chain_762..inv  (.\notGate[761]_keep (notGate_761), 
            .\notGate[762] (notGate_762)) /* synthesis syn_module_defined=1 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(32[13:44])
    inverter_U264 \inverter_chain_761..inv  (.\notGate[760]_keep (notGate_760), 
            .\notGate[761] (notGate_761)) /* synthesis syn_module_defined=1 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(32[13:44])
    inverter_U265 \inverter_chain_760..inv  (.\notGate[759]_keep (notGate_759), 
            .\notGate[760] (notGate_760)) /* synthesis syn_module_defined=1 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(32[13:44])
    inverter_U266 \inverter_chain_75..inv  (.\notGate[74]_keep (notGate_74), 
            .\notGate[75] (notGate_75)) /* synthesis syn_module_defined=1 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(32[13:44])
    inverter_U267 \inverter_chain_759..inv  (.\notGate[758]_keep (notGate_758), 
            .\notGate[759] (notGate_759)) /* synthesis syn_module_defined=1 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(32[13:44])
    inverter_U268 \inverter_chain_758..inv  (.\notGate[757]_keep (notGate_757), 
            .\notGate[758] (notGate_758)) /* synthesis syn_module_defined=1 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(32[13:44])
    inverter_U269 \inverter_chain_757..inv  (.\notGate[756]_keep (notGate_756), 
            .\notGate[757] (notGate_757)) /* synthesis syn_module_defined=1 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(32[13:44])
    inverter_U270 \inverter_chain_756..inv  (.\notGate[755]_keep (notGate_755), 
            .\notGate[756] (notGate_756)) /* synthesis syn_module_defined=1 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(32[13:44])
    inverter_U271 \inverter_chain_755..inv  (.\notGate[754]_keep (notGate_754), 
            .\notGate[755] (notGate_755)) /* synthesis syn_module_defined=1 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(32[13:44])
    inverter_U272 \inverter_chain_754..inv  (.\notGate[753]_keep (notGate_753), 
            .\notGate[754] (notGate_754)) /* synthesis syn_module_defined=1 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(32[13:44])
    inverter_U273 \inverter_chain_753..inv  (.\notGate[752]_keep (notGate_752), 
            .\notGate[753] (notGate_753)) /* synthesis syn_module_defined=1 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(32[13:44])
    inverter_U274 \inverter_chain_752..inv  (.\notGate[751]_keep (notGate_751), 
            .\notGate[752] (notGate_752)) /* synthesis syn_module_defined=1 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(32[13:44])
    inverter_U275 \inverter_chain_751..inv  (.\notGate[750]_keep (notGate_750), 
            .\notGate[751] (notGate_751)) /* synthesis syn_module_defined=1 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(32[13:44])
    inverter_U276 \inverter_chain_750..inv  (.\notGate[749]_keep (notGate_749), 
            .\notGate[750] (notGate_750)) /* synthesis syn_module_defined=1 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(32[13:44])
    inverter_U277 \inverter_chain_74..inv  (.\notGate[73]_keep (notGate_73), 
            .\notGate[74] (notGate_74)) /* synthesis syn_module_defined=1 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(32[13:44])
    inverter_U278 \inverter_chain_749..inv  (.\notGate[748]_keep (notGate_748), 
            .\notGate[749] (notGate_749)) /* synthesis syn_module_defined=1 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(32[13:44])
    inverter_U279 \inverter_chain_748..inv  (.\notGate[747]_keep (notGate_747), 
            .\notGate[748] (notGate_748)) /* synthesis syn_module_defined=1 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(32[13:44])
    inverter_U280 \inverter_chain_747..inv  (.\notGate[746]_keep (notGate_746), 
            .\notGate[747] (notGate_747)) /* synthesis syn_module_defined=1 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(32[13:44])
    inverter_U281 \inverter_chain_746..inv  (.\notGate[745]_keep (notGate_745), 
            .\notGate[746] (notGate_746)) /* synthesis syn_module_defined=1 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(32[13:44])
    inverter_U282 \inverter_chain_745..inv  (.\notGate[744]_keep (notGate_744), 
            .\notGate[745] (notGate_745)) /* synthesis syn_module_defined=1 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(32[13:44])
    inverter_U283 \inverter_chain_744..inv  (.\notGate[743]_keep (notGate_743), 
            .\notGate[744] (notGate_744)) /* synthesis syn_module_defined=1 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(32[13:44])
    inverter_U284 \inverter_chain_743..inv  (.\notGate[742]_keep (notGate_742), 
            .\notGate[743] (notGate_743)) /* synthesis syn_module_defined=1 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(32[13:44])
    inverter_U285 \inverter_chain_742..inv  (.\notGate[741]_keep (notGate_741), 
            .\notGate[742] (notGate_742)) /* synthesis syn_module_defined=1 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(32[13:44])
    inverter_U286 \inverter_chain_741..inv  (.\notGate[740]_keep (notGate_740), 
            .\notGate[741] (notGate_741)) /* synthesis syn_module_defined=1 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(32[13:44])
    inverter_U287 \inverter_chain_740..inv  (.\notGate[739]_keep (notGate_739), 
            .\notGate[740] (notGate_740)) /* synthesis syn_module_defined=1 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(32[13:44])
    inverter_U288 \inverter_chain_73..inv  (.\notGate[72]_keep (notGate_72), 
            .\notGate[73] (notGate_73)) /* synthesis syn_module_defined=1 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(32[13:44])
    inverter_U289 \inverter_chain_739..inv  (.\notGate[738]_keep (notGate_738), 
            .\notGate[739] (notGate_739)) /* synthesis syn_module_defined=1 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(32[13:44])
    inverter_U290 \inverter_chain_738..inv  (.\notGate[737]_keep (notGate_737), 
            .\notGate[738] (notGate_738)) /* synthesis syn_module_defined=1 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(32[13:44])
    inverter_U291 \inverter_chain_737..inv  (.\notGate[736]_keep (notGate_736), 
            .\notGate[737] (notGate_737)) /* synthesis syn_module_defined=1 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(32[13:44])
    inverter_U292 \inverter_chain_736..inv  (.\notGate[735]_keep (notGate_735), 
            .\notGate[736] (notGate_736)) /* synthesis syn_module_defined=1 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(32[13:44])
    inverter_U293 \inverter_chain_735..inv  (.\notGate[734]_keep (notGate_734), 
            .\notGate[735] (notGate_735)) /* synthesis syn_module_defined=1 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(32[13:44])
    inverter_U294 \inverter_chain_734..inv  (.\notGate[733]_keep (notGate_733), 
            .\notGate[734] (notGate_734)) /* synthesis syn_module_defined=1 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(32[13:44])
    inverter_U295 \inverter_chain_733..inv  (.\notGate[732]_keep (notGate_732), 
            .\notGate[733] (notGate_733)) /* synthesis syn_module_defined=1 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(32[13:44])
    inverter_U296 \inverter_chain_732..inv  (.\notGate[731]_keep (notGate_731), 
            .\notGate[732] (notGate_732)) /* synthesis syn_module_defined=1 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(32[13:44])
    inverter_U297 \inverter_chain_731..inv  (.\notGate[730]_keep (notGate_730), 
            .\notGate[731] (notGate_731)) /* synthesis syn_module_defined=1 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(32[13:44])
    inverter_U298 \inverter_chain_730..inv  (.\notGate[729]_keep (notGate_729), 
            .\notGate[730] (notGate_730)) /* synthesis syn_module_defined=1 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(32[13:44])
    inverter_U299 \inverter_chain_72..inv  (.\notGate[71]_keep (notGate_71), 
            .\notGate[72] (notGate_72)) /* synthesis syn_module_defined=1 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(32[13:44])
    inverter_U300 \inverter_chain_729..inv  (.\notGate[728]_keep (notGate_728), 
            .\notGate[729] (notGate_729)) /* synthesis syn_module_defined=1 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(32[13:44])
    inverter_U301 \inverter_chain_728..inv  (.\notGate[727]_keep (notGate_727), 
            .\notGate[728] (notGate_728)) /* synthesis syn_module_defined=1 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(32[13:44])
    inverter_U302 \inverter_chain_727..inv  (.\notGate[726]_keep (notGate_726), 
            .\notGate[727] (notGate_727)) /* synthesis syn_module_defined=1 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(32[13:44])
    inverter_U303 \inverter_chain_726..inv  (.\notGate[725]_keep (notGate_725), 
            .\notGate[726] (notGate_726)) /* synthesis syn_module_defined=1 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(32[13:44])
    inverter_U304 \inverter_chain_725..inv  (.\notGate[724]_keep (notGate_724), 
            .\notGate[725] (notGate_725)) /* synthesis syn_module_defined=1 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(32[13:44])
    inverter_U305 \inverter_chain_724..inv  (.\notGate[723]_keep (notGate_723), 
            .\notGate[724] (notGate_724)) /* synthesis syn_module_defined=1 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(32[13:44])
    inverter_U306 \inverter_chain_723..inv  (.\notGate[722]_keep (notGate_722), 
            .\notGate[723] (notGate_723)) /* synthesis syn_module_defined=1 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(32[13:44])
    inverter_U307 \inverter_chain_722..inv  (.\notGate[721]_keep (notGate_721), 
            .\notGate[722] (notGate_722)) /* synthesis syn_module_defined=1 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(32[13:44])
    inverter_U308 \inverter_chain_721..inv  (.\notGate[720]_keep (notGate_720), 
            .\notGate[721] (notGate_721)) /* synthesis syn_module_defined=1 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(32[13:44])
    inverter_U309 \inverter_chain_720..inv  (.\notGate[719]_keep (notGate_719), 
            .\notGate[720] (notGate_720)) /* synthesis syn_module_defined=1 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(32[13:44])
    inverter_U310 \inverter_chain_71..inv  (.\notGate[70]_keep (notGate_70), 
            .\notGate[71] (notGate_71)) /* synthesis syn_module_defined=1 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(32[13:44])
    inverter_U311 \inverter_chain_719..inv  (.\notGate[718]_keep (notGate_718), 
            .\notGate[719] (notGate_719)) /* synthesis syn_module_defined=1 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(32[13:44])
    inverter_U312 \inverter_chain_718..inv  (.\notGate[717]_keep (notGate_717), 
            .\notGate[718] (notGate_718)) /* synthesis syn_module_defined=1 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(32[13:44])
    inverter_U313 \inverter_chain_717..inv  (.\notGate[716]_keep (notGate_716), 
            .\notGate[717] (notGate_717)) /* synthesis syn_module_defined=1 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(32[13:44])
    inverter_U314 \inverter_chain_716..inv  (.\notGate[715]_keep (notGate_715), 
            .\notGate[716] (notGate_716)) /* synthesis syn_module_defined=1 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(32[13:44])
    inverter_U315 \inverter_chain_715..inv  (.\notGate[714]_keep (notGate_714), 
            .\notGate[715] (notGate_715)) /* synthesis syn_module_defined=1 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(32[13:44])
    inverter_U316 \inverter_chain_714..inv  (.\notGate[713]_keep (notGate_713), 
            .\notGate[714] (notGate_714)) /* synthesis syn_module_defined=1 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(32[13:44])
    inverter_U317 \inverter_chain_713..inv  (.\notGate[712]_keep (notGate_712), 
            .\notGate[713] (notGate_713)) /* synthesis syn_module_defined=1 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(32[13:44])
    inverter_U318 \inverter_chain_712..inv  (.\notGate[711]_keep (notGate_711), 
            .\notGate[712] (notGate_712)) /* synthesis syn_module_defined=1 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(32[13:44])
    inverter_U319 \inverter_chain_711..inv  (.\notGate[710]_keep (notGate_710), 
            .\notGate[711] (notGate_711)) /* synthesis syn_module_defined=1 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(32[13:44])
    inverter_U320 \inverter_chain_710..inv  (.\notGate[709]_keep (notGate_709), 
            .\notGate[710] (notGate_710)) /* synthesis syn_module_defined=1 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(32[13:44])
    inverter_U321 \inverter_chain_70..inv  (.\notGate[69]_keep (notGate_69), 
            .\notGate[70] (notGate_70)) /* synthesis syn_module_defined=1 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(32[13:44])
    inverter_U322 \inverter_chain_709..inv  (.\notGate[708]_keep (notGate_708), 
            .\notGate[709] (notGate_709)) /* synthesis syn_module_defined=1 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(32[13:44])
    inverter_U323 \inverter_chain_708..inv  (.\notGate[707]_keep (notGate_707), 
            .\notGate[708] (notGate_708)) /* synthesis syn_module_defined=1 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(32[13:44])
    inverter_U324 \inverter_chain_707..inv  (.\notGate[706]_keep (notGate_706), 
            .\notGate[707] (notGate_707)) /* synthesis syn_module_defined=1 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(32[13:44])
    inverter_U325 \inverter_chain_706..inv  (.\notGate[705]_keep (notGate_705), 
            .\notGate[706] (notGate_706)) /* synthesis syn_module_defined=1 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(32[13:44])
    inverter_U326 \inverter_chain_705..inv  (.\notGate[704]_keep (notGate_704), 
            .\notGate[705] (notGate_705)) /* synthesis syn_module_defined=1 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(32[13:44])
    inverter_U327 \inverter_chain_704..inv  (.\notGate[703]_keep (notGate_703), 
            .\notGate[704] (notGate_704)) /* synthesis syn_module_defined=1 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(32[13:44])
    inverter_U328 \inverter_chain_703..inv  (.\notGate[702]_keep (notGate_702), 
            .\notGate[703] (notGate_703)) /* synthesis syn_module_defined=1 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(32[13:44])
    inverter_U329 \inverter_chain_702..inv  (.\notGate[701]_keep (notGate_701), 
            .\notGate[702] (notGate_702)) /* synthesis syn_module_defined=1 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(32[13:44])
    inverter_U330 \inverter_chain_701..inv  (.\notGate[700]_keep (notGate_700), 
            .\notGate[701] (notGate_701)) /* synthesis syn_module_defined=1 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(32[13:44])
    inverter_U331 \inverter_chain_700..inv  (.\notGate[699]_keep (notGate_699), 
            .\notGate[700] (notGate_700)) /* synthesis syn_module_defined=1 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(32[13:44])
    inverter_U332 \inverter_chain_6..inv  (.\notGate[5]_keep (notGate_5), 
            .\notGate[6] (notGate_6)) /* synthesis syn_module_defined=1 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(32[13:44])
    inverter_U333 \inverter_chain_69..inv  (.\notGate[68]_keep (notGate_68), 
            .\notGate[69] (notGate_69)) /* synthesis syn_module_defined=1 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(32[13:44])
    inverter_U334 \inverter_chain_699..inv  (.\notGate[698]_keep (notGate_698), 
            .\notGate[699] (notGate_699)) /* synthesis syn_module_defined=1 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(32[13:44])
    inverter_U335 \inverter_chain_698..inv  (.\notGate[697]_keep (notGate_697), 
            .\notGate[698] (notGate_698)) /* synthesis syn_module_defined=1 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(32[13:44])
    inverter_U336 \inverter_chain_697..inv  (.\notGate[696]_keep (notGate_696), 
            .\notGate[697] (notGate_697)) /* synthesis syn_module_defined=1 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(32[13:44])
    inverter_U337 \inverter_chain_696..inv  (.\notGate[695]_keep (notGate_695), 
            .\notGate[696] (notGate_696)) /* synthesis syn_module_defined=1 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(32[13:44])
    inverter_U338 \inverter_chain_695..inv  (.\notGate[694]_keep (notGate_694), 
            .\notGate[695] (notGate_695)) /* synthesis syn_module_defined=1 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(32[13:44])
    inverter_U339 \inverter_chain_694..inv  (.\notGate[693]_keep (notGate_693), 
            .\notGate[694] (notGate_694)) /* synthesis syn_module_defined=1 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(32[13:44])
    inverter_U340 \inverter_chain_693..inv  (.\notGate[692]_keep (notGate_692), 
            .\notGate[693] (notGate_693)) /* synthesis syn_module_defined=1 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(32[13:44])
    inverter_U341 \inverter_chain_692..inv  (.\notGate[691]_keep (notGate_691), 
            .\notGate[692] (notGate_692)) /* synthesis syn_module_defined=1 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(32[13:44])
    inverter_U342 \inverter_chain_691..inv  (.\notGate[690]_keep (notGate_690), 
            .\notGate[691] (notGate_691)) /* synthesis syn_module_defined=1 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(32[13:44])
    inverter_U343 \inverter_chain_690..inv  (.\notGate[689]_keep (notGate_689), 
            .\notGate[690] (notGate_690)) /* synthesis syn_module_defined=1 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(32[13:44])
    inverter_U344 \inverter_chain_68..inv  (.\notGate[67]_keep (notGate_67), 
            .\notGate[68] (notGate_68)) /* synthesis syn_module_defined=1 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(32[13:44])
    inverter_U345 \inverter_chain_689..inv  (.\notGate[688]_keep (notGate_688), 
            .\notGate[689] (notGate_689)) /* synthesis syn_module_defined=1 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(32[13:44])
    inverter_U346 \inverter_chain_688..inv  (.\notGate[687]_keep (notGate_687), 
            .\notGate[688] (notGate_688)) /* synthesis syn_module_defined=1 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(32[13:44])
    inverter_U347 \inverter_chain_687..inv  (.\notGate[686]_keep (notGate_686), 
            .\notGate[687] (notGate_687)) /* synthesis syn_module_defined=1 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(32[13:44])
    inverter_U348 \inverter_chain_686..inv  (.\notGate[685]_keep (notGate_685), 
            .\notGate[686] (notGate_686)) /* synthesis syn_module_defined=1 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(32[13:44])
    inverter_U349 \inverter_chain_685..inv  (.\notGate[684]_keep (notGate_684), 
            .\notGate[685] (notGate_685)) /* synthesis syn_module_defined=1 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(32[13:44])
    inverter_U350 \inverter_chain_684..inv  (.\notGate[683]_keep (notGate_683), 
            .\notGate[684] (notGate_684)) /* synthesis syn_module_defined=1 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(32[13:44])
    inverter_U351 \inverter_chain_683..inv  (.\notGate[682]_keep (notGate_682), 
            .\notGate[683] (notGate_683)) /* synthesis syn_module_defined=1 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(32[13:44])
    inverter_U352 \inverter_chain_682..inv  (.\notGate[681]_keep (notGate_681), 
            .\notGate[682] (notGate_682)) /* synthesis syn_module_defined=1 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(32[13:44])
    inverter_U353 \inverter_chain_681..inv  (.\notGate[680]_keep (notGate_680), 
            .\notGate[681] (notGate_681)) /* synthesis syn_module_defined=1 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(32[13:44])
    inverter_U354 \inverter_chain_680..inv  (.\notGate[679]_keep (notGate_679), 
            .\notGate[680] (notGate_680)) /* synthesis syn_module_defined=1 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(32[13:44])
    inverter_U355 \inverter_chain_67..inv  (.\notGate[66]_keep (notGate_66), 
            .\notGate[67] (notGate_67)) /* synthesis syn_module_defined=1 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(32[13:44])
    inverter_U356 \inverter_chain_679..inv  (.\notGate[678]_keep (notGate_678), 
            .\notGate[679] (notGate_679)) /* synthesis syn_module_defined=1 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(32[13:44])
    inverter_U357 \inverter_chain_678..inv  (.\notGate[677]_keep (notGate_677), 
            .\notGate[678] (notGate_678)) /* synthesis syn_module_defined=1 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(32[13:44])
    inverter_U358 \inverter_chain_677..inv  (.\notGate[676]_keep (notGate_676), 
            .\notGate[677] (notGate_677)) /* synthesis syn_module_defined=1 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(32[13:44])
    inverter_U359 \inverter_chain_676..inv  (.\notGate[675]_keep (notGate_675), 
            .\notGate[676] (notGate_676)) /* synthesis syn_module_defined=1 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(32[13:44])
    inverter_U360 \inverter_chain_675..inv  (.\notGate[674]_keep (notGate_674), 
            .\notGate[675] (notGate_675)) /* synthesis syn_module_defined=1 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(32[13:44])
    inverter_U361 \inverter_chain_674..inv  (.\notGate[673]_keep (notGate_673), 
            .\notGate[674] (notGate_674)) /* synthesis syn_module_defined=1 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(32[13:44])
    inverter_U362 \inverter_chain_673..inv  (.\notGate[672]_keep (notGate_672), 
            .\notGate[673] (notGate_673)) /* synthesis syn_module_defined=1 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(32[13:44])
    inverter_U363 \inverter_chain_672..inv  (.\notGate[671]_keep (notGate_671), 
            .\notGate[672] (notGate_672)) /* synthesis syn_module_defined=1 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(32[13:44])
    inverter_U364 \inverter_chain_671..inv  (.\notGate[670]_keep (notGate_670), 
            .\notGate[671] (notGate_671)) /* synthesis syn_module_defined=1 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(32[13:44])
    inverter_U365 \inverter_chain_670..inv  (.\notGate[669]_keep (notGate_669), 
            .\notGate[670] (notGate_670)) /* synthesis syn_module_defined=1 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(32[13:44])
    inverter_U366 \inverter_chain_66..inv  (.\notGate[65]_keep (notGate_65), 
            .\notGate[66] (notGate_66)) /* synthesis syn_module_defined=1 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(32[13:44])
    inverter_U367 \inverter_chain_669..inv  (.\notGate[668]_keep (notGate_668), 
            .\notGate[669] (notGate_669)) /* synthesis syn_module_defined=1 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(32[13:44])
    inverter_U368 \inverter_chain_668..inv  (.\notGate[667]_keep (notGate_667), 
            .\notGate[668] (notGate_668)) /* synthesis syn_module_defined=1 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(32[13:44])
    inverter_U369 \inverter_chain_667..inv  (.\notGate[666]_keep (notGate_666), 
            .\notGate[667] (notGate_667)) /* synthesis syn_module_defined=1 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(32[13:44])
    inverter_U370 \inverter_chain_666..inv  (.\notGate[665]_keep (notGate_665), 
            .\notGate[666] (notGate_666)) /* synthesis syn_module_defined=1 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(32[13:44])
    inverter_U371 \inverter_chain_665..inv  (.\notGate[664]_keep (notGate_664), 
            .\notGate[665] (notGate_665)) /* synthesis syn_module_defined=1 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(32[13:44])
    inverter_U372 \inverter_chain_664..inv  (.\notGate[663]_keep (notGate_663), 
            .\notGate[664] (notGate_664)) /* synthesis syn_module_defined=1 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(32[13:44])
    inverter_U373 \inverter_chain_663..inv  (.\notGate[662]_keep (notGate_662), 
            .\notGate[663] (notGate_663)) /* synthesis syn_module_defined=1 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(32[13:44])
    inverter_U374 \inverter_chain_662..inv  (.\notGate[661]_keep (notGate_661), 
            .\notGate[662] (notGate_662)) /* synthesis syn_module_defined=1 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(32[13:44])
    inverter_U375 \inverter_chain_661..inv  (.\notGate[660]_keep (notGate_660), 
            .\notGate[661] (notGate_661)) /* synthesis syn_module_defined=1 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(32[13:44])
    inverter_U376 \inverter_chain_660..inv  (.\notGate[659]_keep (notGate_659), 
            .\notGate[660] (notGate_660)) /* synthesis syn_module_defined=1 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(32[13:44])
    inverter_U377 \inverter_chain_65..inv  (.\notGate[64]_keep (notGate_64), 
            .\notGate[65] (notGate_65)) /* synthesis syn_module_defined=1 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(32[13:44])
    inverter_U378 \inverter_chain_659..inv  (.\notGate[658]_keep (notGate_658), 
            .\notGate[659] (notGate_659)) /* synthesis syn_module_defined=1 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(32[13:44])
    inverter_U379 \inverter_chain_658..inv  (.\notGate[657]_keep (notGate_657), 
            .\notGate[658] (notGate_658)) /* synthesis syn_module_defined=1 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(32[13:44])
    inverter_U380 \inverter_chain_657..inv  (.\notGate[656]_keep (notGate_656), 
            .\notGate[657] (notGate_657)) /* synthesis syn_module_defined=1 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(32[13:44])
    inverter_U381 \inverter_chain_656..inv  (.\notGate[655]_keep (notGate_655), 
            .\notGate[656] (notGate_656)) /* synthesis syn_module_defined=1 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(32[13:44])
    inverter_U382 \inverter_chain_655..inv  (.\notGate[654]_keep (notGate_654), 
            .\notGate[655] (notGate_655)) /* synthesis syn_module_defined=1 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(32[13:44])
    inverter_U383 \inverter_chain_654..inv  (.\notGate[653]_keep (notGate_653), 
            .\notGate[654] (notGate_654)) /* synthesis syn_module_defined=1 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(32[13:44])
    inverter_U384 \inverter_chain_653..inv  (.\notGate[652]_keep (notGate_652), 
            .\notGate[653] (notGate_653)) /* synthesis syn_module_defined=1 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(32[13:44])
    inverter_U385 \inverter_chain_652..inv  (.\notGate[651]_keep (notGate_651), 
            .\notGate[652] (notGate_652)) /* synthesis syn_module_defined=1 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(32[13:44])
    inverter_U386 \inverter_chain_651..inv  (.\notGate[650]_keep (notGate_650), 
            .\notGate[651] (notGate_651)) /* synthesis syn_module_defined=1 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(32[13:44])
    inverter_U387 \inverter_chain_650..inv  (.\notGate[649]_keep (notGate_649), 
            .\notGate[650] (notGate_650)) /* synthesis syn_module_defined=1 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(32[13:44])
    inverter_U388 \inverter_chain_64..inv  (.\notGate[63]_keep (notGate_63), 
            .\notGate[64] (notGate_64)) /* synthesis syn_module_defined=1 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(32[13:44])
    inverter_U389 \inverter_chain_649..inv  (.\notGate[648]_keep (notGate_648), 
            .\notGate[649] (notGate_649)) /* synthesis syn_module_defined=1 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(32[13:44])
    inverter_U390 \inverter_chain_648..inv  (.\notGate[647]_keep (notGate_647), 
            .\notGate[648] (notGate_648)) /* synthesis syn_module_defined=1 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(32[13:44])
    inverter_U391 \inverter_chain_647..inv  (.\notGate[646]_keep (notGate_646), 
            .\notGate[647] (notGate_647)) /* synthesis syn_module_defined=1 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(32[13:44])
    inverter_U392 \inverter_chain_646..inv  (.\notGate[645]_keep (notGate_645), 
            .\notGate[646] (notGate_646)) /* synthesis syn_module_defined=1 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(32[13:44])
    inverter_U393 \inverter_chain_645..inv  (.\notGate[644]_keep (notGate_644), 
            .\notGate[645] (notGate_645)) /* synthesis syn_module_defined=1 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(32[13:44])
    inverter_U394 \inverter_chain_644..inv  (.\notGate[643]_keep (notGate_643), 
            .\notGate[644] (notGate_644)) /* synthesis syn_module_defined=1 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(32[13:44])
    inverter_U395 \inverter_chain_643..inv  (.\notGate[642]_keep (notGate_642), 
            .\notGate[643] (notGate_643)) /* synthesis syn_module_defined=1 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(32[13:44])
    inverter_U396 \inverter_chain_642..inv  (.\notGate[641]_keep (notGate_641), 
            .\notGate[642] (notGate_642)) /* synthesis syn_module_defined=1 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(32[13:44])
    inverter_U397 \inverter_chain_641..inv  (.\notGate[640]_keep (notGate_640), 
            .\notGate[641] (notGate_641)) /* synthesis syn_module_defined=1 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(32[13:44])
    inverter_U398 \inverter_chain_640..inv  (.\notGate[639]_keep (notGate_639), 
            .\notGate[640] (notGate_640)) /* synthesis syn_module_defined=1 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(32[13:44])
    inverter_U399 \inverter_chain_63..inv  (.\notGate[62]_keep (notGate_62), 
            .\notGate[63] (notGate_63)) /* synthesis syn_module_defined=1 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(32[13:44])
    inverter_U400 \inverter_chain_639..inv  (.\notGate[638]_keep (notGate_638), 
            .\notGate[639] (notGate_639)) /* synthesis syn_module_defined=1 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(32[13:44])
    inverter_U401 \inverter_chain_638..inv  (.\notGate[637]_keep (notGate_637), 
            .\notGate[638] (notGate_638)) /* synthesis syn_module_defined=1 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(32[13:44])
    inverter_U402 \inverter_chain_637..inv  (.\notGate[636]_keep (notGate_636), 
            .\notGate[637] (notGate_637)) /* synthesis syn_module_defined=1 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(32[13:44])
    inverter_U403 \inverter_chain_636..inv  (.\notGate[635]_keep (notGate_635), 
            .\notGate[636] (notGate_636)) /* synthesis syn_module_defined=1 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(32[13:44])
    inverter_U404 \inverter_chain_635..inv  (.\notGate[634]_keep (notGate_634), 
            .\notGate[635] (notGate_635)) /* synthesis syn_module_defined=1 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(32[13:44])
    inverter_U405 \inverter_chain_634..inv  (.\notGate[633]_keep (notGate_633), 
            .\notGate[634] (notGate_634)) /* synthesis syn_module_defined=1 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(32[13:44])
    inverter_U406 \inverter_chain_633..inv  (.\notGate[632]_keep (notGate_632), 
            .\notGate[633] (notGate_633)) /* synthesis syn_module_defined=1 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(32[13:44])
    inverter_U407 \inverter_chain_632..inv  (.\notGate[631]_keep (notGate_631), 
            .\notGate[632] (notGate_632)) /* synthesis syn_module_defined=1 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(32[13:44])
    inverter_U408 \inverter_chain_631..inv  (.\notGate[630]_keep (notGate_630), 
            .\notGate[631] (notGate_631)) /* synthesis syn_module_defined=1 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(32[13:44])
    inverter_U409 \inverter_chain_630..inv  (.\notGate[629]_keep (notGate_629), 
            .\notGate[630] (notGate_630)) /* synthesis syn_module_defined=1 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(32[13:44])
    inverter_U410 \inverter_chain_62..inv  (.\notGate[61]_keep (notGate_61), 
            .\notGate[62] (notGate_62)) /* synthesis syn_module_defined=1 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(32[13:44])
    inverter_U411 \inverter_chain_629..inv  (.\notGate[628]_keep (notGate_628), 
            .\notGate[629] (notGate_629)) /* synthesis syn_module_defined=1 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(32[13:44])
    inverter_U412 \inverter_chain_628..inv  (.\notGate[627]_keep (notGate_627), 
            .\notGate[628] (notGate_628)) /* synthesis syn_module_defined=1 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(32[13:44])
    inverter_U413 \inverter_chain_627..inv  (.\notGate[626]_keep (notGate_626), 
            .\notGate[627] (notGate_627)) /* synthesis syn_module_defined=1 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(32[13:44])
    inverter_U414 \inverter_chain_626..inv  (.\notGate[625]_keep (notGate_625), 
            .\notGate[626] (notGate_626)) /* synthesis syn_module_defined=1 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(32[13:44])
    inverter_U415 \inverter_chain_625..inv  (.\notGate[624]_keep (notGate_624), 
            .\notGate[625] (notGate_625)) /* synthesis syn_module_defined=1 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(32[13:44])
    inverter_U416 \inverter_chain_624..inv  (.\notGate[623]_keep (notGate_623), 
            .\notGate[624] (notGate_624)) /* synthesis syn_module_defined=1 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(32[13:44])
    inverter_U417 \inverter_chain_623..inv  (.\notGate[622]_keep (notGate_622), 
            .\notGate[623] (notGate_623)) /* synthesis syn_module_defined=1 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(32[13:44])
    inverter_U418 \inverter_chain_622..inv  (.\notGate[621]_keep (notGate_621), 
            .\notGate[622] (notGate_622)) /* synthesis syn_module_defined=1 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(32[13:44])
    inverter_U419 \inverter_chain_621..inv  (.\notGate[620]_keep (notGate_620), 
            .\notGate[621] (notGate_621)) /* synthesis syn_module_defined=1 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(32[13:44])
    inverter_U420 \inverter_chain_620..inv  (.\notGate[619]_keep (notGate_619), 
            .\notGate[620] (notGate_620)) /* synthesis syn_module_defined=1 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(32[13:44])
    inverter_U421 \inverter_chain_61..inv  (.\notGate[60]_keep (notGate_60), 
            .\notGate[61] (notGate_61)) /* synthesis syn_module_defined=1 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(32[13:44])
    inverter_U422 \inverter_chain_619..inv  (.\notGate[618]_keep (notGate_618), 
            .\notGate[619] (notGate_619)) /* synthesis syn_module_defined=1 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(32[13:44])
    inverter_U423 \inverter_chain_618..inv  (.\notGate[617]_keep (notGate_617), 
            .\notGate[618] (notGate_618)) /* synthesis syn_module_defined=1 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(32[13:44])
    inverter_U424 \inverter_chain_617..inv  (.\notGate[616]_keep (notGate_616), 
            .\notGate[617] (notGate_617)) /* synthesis syn_module_defined=1 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(32[13:44])
    inverter_U425 \inverter_chain_616..inv  (.\notGate[615]_keep (notGate_615), 
            .\notGate[616] (notGate_616)) /* synthesis syn_module_defined=1 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(32[13:44])
    inverter_U426 \inverter_chain_615..inv  (.\notGate[614]_keep (notGate_614), 
            .\notGate[615] (notGate_615)) /* synthesis syn_module_defined=1 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(32[13:44])
    inverter_U427 \inverter_chain_614..inv  (.\notGate[613]_keep (notGate_613), 
            .\notGate[614] (notGate_614)) /* synthesis syn_module_defined=1 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(32[13:44])
    inverter_U428 \inverter_chain_613..inv  (.\notGate[612]_keep (notGate_612), 
            .\notGate[613] (notGate_613)) /* synthesis syn_module_defined=1 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(32[13:44])
    inverter_U429 \inverter_chain_612..inv  (.\notGate[611]_keep (notGate_611), 
            .\notGate[612] (notGate_612)) /* synthesis syn_module_defined=1 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(32[13:44])
    inverter_U430 \inverter_chain_611..inv  (.\notGate[610]_keep (notGate_610), 
            .\notGate[611] (notGate_611)) /* synthesis syn_module_defined=1 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(32[13:44])
    inverter_U431 \inverter_chain_610..inv  (.\notGate[609]_keep (notGate_609), 
            .\notGate[610] (notGate_610)) /* synthesis syn_module_defined=1 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(32[13:44])
    inverter_U432 \inverter_chain_60..inv  (.\notGate[59]_keep (notGate_59), 
            .\notGate[60] (notGate_60)) /* synthesis syn_module_defined=1 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(32[13:44])
    inverter_U433 \inverter_chain_609..inv  (.\notGate[608]_keep (notGate_608), 
            .\notGate[609] (notGate_609)) /* synthesis syn_module_defined=1 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(32[13:44])
    inverter_U434 \inverter_chain_608..inv  (.\notGate[607]_keep (notGate_607), 
            .\notGate[608] (notGate_608)) /* synthesis syn_module_defined=1 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(32[13:44])
    inverter_U435 \inverter_chain_607..inv  (.\notGate[606]_keep (notGate_606), 
            .\notGate[607] (notGate_607)) /* synthesis syn_module_defined=1 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(32[13:44])
    inverter_U436 \inverter_chain_606..inv  (.\notGate[605]_keep (notGate_605), 
            .\notGate[606] (notGate_606)) /* synthesis syn_module_defined=1 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(32[13:44])
    inverter_U437 \inverter_chain_605..inv  (.\notGate[604]_keep (notGate_604), 
            .\notGate[605] (notGate_605)) /* synthesis syn_module_defined=1 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(32[13:44])
    inverter_U438 \inverter_chain_604..inv  (.\notGate[603]_keep (notGate_603), 
            .\notGate[604] (notGate_604)) /* synthesis syn_module_defined=1 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(32[13:44])
    inverter_U439 \inverter_chain_603..inv  (.\notGate[602]_keep (notGate_602), 
            .\notGate[603] (notGate_603)) /* synthesis syn_module_defined=1 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(32[13:44])
    inverter_U440 \inverter_chain_602..inv  (.\notGate[601]_keep (notGate_601), 
            .\notGate[602] (notGate_602)) /* synthesis syn_module_defined=1 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(32[13:44])
    inverter_U441 \inverter_chain_601..inv  (.\notGate[600]_keep (notGate_600), 
            .\notGate[601] (notGate_601)) /* synthesis syn_module_defined=1 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(32[13:44])
    inverter_U442 \inverter_chain_600..inv  (.\notGate[599]_keep (notGate_599), 
            .\notGate[600] (notGate_600)) /* synthesis syn_module_defined=1 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(32[13:44])
    inverter_U443 \inverter_chain_5..inv  (.\notGate[4]_keep (notGate_4), 
            .\notGate[5] (notGate_5)) /* synthesis syn_module_defined=1 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(32[13:44])
    inverter_U444 \inverter_chain_59..inv  (.\notGate[58]_keep (notGate_58), 
            .\notGate[59] (notGate_59)) /* synthesis syn_module_defined=1 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(32[13:44])
    inverter_U445 \inverter_chain_599..inv  (.\notGate[598]_keep (notGate_598), 
            .\notGate[599] (notGate_599)) /* synthesis syn_module_defined=1 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(32[13:44])
    inverter_U446 \inverter_chain_598..inv  (.\notGate[597]_keep (notGate_597), 
            .\notGate[598] (notGate_598)) /* synthesis syn_module_defined=1 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(32[13:44])
    inverter_U447 \inverter_chain_597..inv  (.\notGate[596]_keep (notGate_596), 
            .\notGate[597] (notGate_597)) /* synthesis syn_module_defined=1 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(32[13:44])
    inverter_U448 \inverter_chain_596..inv  (.\notGate[595]_keep (notGate_595), 
            .\notGate[596] (notGate_596)) /* synthesis syn_module_defined=1 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(32[13:44])
    inverter_U449 \inverter_chain_595..inv  (.\notGate[594]_keep (notGate_594), 
            .\notGate[595] (notGate_595)) /* synthesis syn_module_defined=1 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(32[13:44])
    inverter_U450 \inverter_chain_594..inv  (.\notGate[593]_keep (notGate_593), 
            .\notGate[594] (notGate_594)) /* synthesis syn_module_defined=1 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(32[13:44])
    inverter_U451 \inverter_chain_593..inv  (.\notGate[592]_keep (notGate_592), 
            .\notGate[593] (notGate_593)) /* synthesis syn_module_defined=1 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(32[13:44])
    inverter_U452 \inverter_chain_592..inv  (.\notGate[591]_keep (notGate_591), 
            .\notGate[592] (notGate_592)) /* synthesis syn_module_defined=1 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(32[13:44])
    inverter_U453 \inverter_chain_591..inv  (.\notGate[590]_keep (notGate_590), 
            .\notGate[591] (notGate_591)) /* synthesis syn_module_defined=1 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(32[13:44])
    inverter_U454 \inverter_chain_590..inv  (.\notGate[589]_keep (notGate_589), 
            .\notGate[590] (notGate_590)) /* synthesis syn_module_defined=1 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(32[13:44])
    inverter_U455 \inverter_chain_58..inv  (.\notGate[57]_keep (notGate_57), 
            .\notGate[58] (notGate_58)) /* synthesis syn_module_defined=1 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(32[13:44])
    inverter_U456 \inverter_chain_589..inv  (.\notGate[588]_keep (notGate_588), 
            .\notGate[589] (notGate_589)) /* synthesis syn_module_defined=1 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(32[13:44])
    inverter_U457 \inverter_chain_588..inv  (.\notGate[587]_keep (notGate_587), 
            .\notGate[588] (notGate_588)) /* synthesis syn_module_defined=1 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(32[13:44])
    inverter_U458 \inverter_chain_587..inv  (.\notGate[586]_keep (notGate_586), 
            .\notGate[587] (notGate_587)) /* synthesis syn_module_defined=1 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(32[13:44])
    inverter_U459 \inverter_chain_586..inv  (.\notGate[585]_keep (notGate_585), 
            .\notGate[586] (notGate_586)) /* synthesis syn_module_defined=1 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(32[13:44])
    inverter_U460 \inverter_chain_585..inv  (.\notGate[584]_keep (notGate_584), 
            .\notGate[585] (notGate_585)) /* synthesis syn_module_defined=1 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(32[13:44])
    inverter_U461 \inverter_chain_584..inv  (.\notGate[583]_keep (notGate_583), 
            .\notGate[584] (notGate_584)) /* synthesis syn_module_defined=1 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(32[13:44])
    inverter_U462 \inverter_chain_583..inv  (.\notGate[582]_keep (notGate_582), 
            .\notGate[583] (notGate_583)) /* synthesis syn_module_defined=1 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(32[13:44])
    inverter_U463 \inverter_chain_582..inv  (.\notGate[581]_keep (notGate_581), 
            .\notGate[582] (notGate_582)) /* synthesis syn_module_defined=1 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(32[13:44])
    inverter_U464 \inverter_chain_581..inv  (.\notGate[580]_keep (notGate_580), 
            .\notGate[581] (notGate_581)) /* synthesis syn_module_defined=1 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(32[13:44])
    inverter_U465 \inverter_chain_580..inv  (.\notGate[579]_keep (notGate_579), 
            .\notGate[580] (notGate_580)) /* synthesis syn_module_defined=1 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(32[13:44])
    inverter_U466 \inverter_chain_57..inv  (.\notGate[56]_keep (notGate_56), 
            .\notGate[57] (notGate_57)) /* synthesis syn_module_defined=1 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(32[13:44])
    inverter_U467 \inverter_chain_579..inv  (.\notGate[578]_keep (notGate_578), 
            .\notGate[579] (notGate_579)) /* synthesis syn_module_defined=1 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(32[13:44])
    inverter_U468 \inverter_chain_578..inv  (.\notGate[577]_keep (notGate_577), 
            .\notGate[578] (notGate_578)) /* synthesis syn_module_defined=1 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(32[13:44])
    inverter_U469 \inverter_chain_577..inv  (.\notGate[576]_keep (notGate_576), 
            .\notGate[577] (notGate_577)) /* synthesis syn_module_defined=1 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(32[13:44])
    inverter_U470 \inverter_chain_576..inv  (.\notGate[575]_keep (notGate_575), 
            .\notGate[576] (notGate_576)) /* synthesis syn_module_defined=1 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(32[13:44])
    inverter_U471 \inverter_chain_575..inv  (.\notGate[574]_keep (notGate_574), 
            .\notGate[575] (notGate_575)) /* synthesis syn_module_defined=1 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(32[13:44])
    inverter_U472 \inverter_chain_574..inv  (.\notGate[573]_keep (notGate_573), 
            .\notGate[574] (notGate_574)) /* synthesis syn_module_defined=1 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(32[13:44])
    inverter_U473 \inverter_chain_573..inv  (.\notGate[572]_keep (notGate_572), 
            .\notGate[573] (notGate_573)) /* synthesis syn_module_defined=1 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(32[13:44])
    inverter_U474 \inverter_chain_572..inv  (.\notGate[571]_keep (notGate_571), 
            .\notGate[572] (notGate_572)) /* synthesis syn_module_defined=1 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(32[13:44])
    inverter_U475 \inverter_chain_571..inv  (.\notGate[570]_keep (notGate_570), 
            .\notGate[571] (notGate_571)) /* synthesis syn_module_defined=1 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(32[13:44])
    inverter_U476 \inverter_chain_570..inv  (.\notGate[569]_keep (notGate_569), 
            .\notGate[570] (notGate_570)) /* synthesis syn_module_defined=1 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(32[13:44])
    inverter_U477 \inverter_chain_56..inv  (.\notGate[55]_keep (notGate_55), 
            .\notGate[56] (notGate_56)) /* synthesis syn_module_defined=1 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(32[13:44])
    inverter_U478 \inverter_chain_569..inv  (.\notGate[568]_keep (notGate_568), 
            .\notGate[569] (notGate_569)) /* synthesis syn_module_defined=1 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(32[13:44])
    inverter_U479 \inverter_chain_568..inv  (.\notGate[567]_keep (notGate_567), 
            .\notGate[568] (notGate_568)) /* synthesis syn_module_defined=1 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(32[13:44])
    inverter_U480 \inverter_chain_567..inv  (.\notGate[566]_keep (notGate_566), 
            .\notGate[567] (notGate_567)) /* synthesis syn_module_defined=1 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(32[13:44])
    inverter_U481 \inverter_chain_566..inv  (.\notGate[565]_keep (notGate_565), 
            .\notGate[566] (notGate_566)) /* synthesis syn_module_defined=1 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(32[13:44])
    inverter_U482 \inverter_chain_565..inv  (.\notGate[564]_keep (notGate_564), 
            .\notGate[565] (notGate_565)) /* synthesis syn_module_defined=1 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(32[13:44])
    inverter_U483 \inverter_chain_564..inv  (.\notGate[563]_keep (notGate_563), 
            .\notGate[564] (notGate_564)) /* synthesis syn_module_defined=1 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(32[13:44])
    inverter_U484 \inverter_chain_563..inv  (.\notGate[562]_keep (notGate_562), 
            .\notGate[563] (notGate_563)) /* synthesis syn_module_defined=1 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(32[13:44])
    inverter_U485 \inverter_chain_562..inv  (.\notGate[561]_keep (notGate_561), 
            .\notGate[562] (notGate_562)) /* synthesis syn_module_defined=1 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(32[13:44])
    inverter_U486 \inverter_chain_561..inv  (.\notGate[560]_keep (notGate_560), 
            .\notGate[561] (notGate_561)) /* synthesis syn_module_defined=1 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(32[13:44])
    inverter_U487 \inverter_chain_560..inv  (.\notGate[559]_keep (notGate_559), 
            .\notGate[560] (notGate_560)) /* synthesis syn_module_defined=1 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(32[13:44])
    inverter_U488 \inverter_chain_55..inv  (.\notGate[54]_keep (notGate_54), 
            .\notGate[55] (notGate_55)) /* synthesis syn_module_defined=1 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(32[13:44])
    inverter_U489 \inverter_chain_559..inv  (.\notGate[558]_keep (notGate_558), 
            .\notGate[559] (notGate_559)) /* synthesis syn_module_defined=1 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(32[13:44])
    inverter_U490 \inverter_chain_558..inv  (.\notGate[557]_keep (notGate_557), 
            .\notGate[558] (notGate_558)) /* synthesis syn_module_defined=1 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(32[13:44])
    inverter_U491 \inverter_chain_557..inv  (.\notGate[556]_keep (notGate_556), 
            .\notGate[557] (notGate_557)) /* synthesis syn_module_defined=1 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(32[13:44])
    inverter_U492 \inverter_chain_556..inv  (.\notGate[555]_keep (notGate_555), 
            .\notGate[556] (notGate_556)) /* synthesis syn_module_defined=1 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(32[13:44])
    inverter_U493 \inverter_chain_555..inv  (.\notGate[554]_keep (notGate_554), 
            .\notGate[555] (notGate_555)) /* synthesis syn_module_defined=1 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(32[13:44])
    inverter_U494 \inverter_chain_554..inv  (.\notGate[553]_keep (notGate_553), 
            .\notGate[554] (notGate_554)) /* synthesis syn_module_defined=1 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(32[13:44])
    inverter_U495 \inverter_chain_553..inv  (.\notGate[552]_keep (notGate_552), 
            .\notGate[553] (notGate_553)) /* synthesis syn_module_defined=1 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(32[13:44])
    inverter_U496 \inverter_chain_552..inv  (.\notGate[551]_keep (notGate_551), 
            .\notGate[552] (notGate_552)) /* synthesis syn_module_defined=1 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(32[13:44])
    inverter_U497 \inverter_chain_551..inv  (.\notGate[550]_keep (notGate_550), 
            .\notGate[551] (notGate_551)) /* synthesis syn_module_defined=1 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(32[13:44])
    inverter_U498 \inverter_chain_550..inv  (.\notGate[549]_keep (notGate_549), 
            .\notGate[550] (notGate_550)) /* synthesis syn_module_defined=1 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(32[13:44])
    inverter_U499 \inverter_chain_54..inv  (.\notGate[53]_keep (notGate_53), 
            .\notGate[54] (notGate_54)) /* synthesis syn_module_defined=1 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(32[13:44])
    inverter_U500 \inverter_chain_549..inv  (.\notGate[548]_keep (notGate_548), 
            .\notGate[549] (notGate_549)) /* synthesis syn_module_defined=1 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(32[13:44])
    inverter_U501 \inverter_chain_548..inv  (.\notGate[547]_keep (notGate_547), 
            .\notGate[548] (notGate_548)) /* synthesis syn_module_defined=1 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(32[13:44])
    inverter_U502 \inverter_chain_547..inv  (.\notGate[546]_keep (notGate_546), 
            .\notGate[547] (notGate_547)) /* synthesis syn_module_defined=1 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(32[13:44])
    inverter_U503 \inverter_chain_546..inv  (.\notGate[545]_keep (notGate_545), 
            .\notGate[546] (notGate_546)) /* synthesis syn_module_defined=1 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(32[13:44])
    inverter_U504 \inverter_chain_545..inv  (.\notGate[544]_keep (notGate_544), 
            .\notGate[545] (notGate_545)) /* synthesis syn_module_defined=1 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(32[13:44])
    inverter_U505 \inverter_chain_544..inv  (.\notGate[543]_keep (notGate_543), 
            .\notGate[544] (notGate_544)) /* synthesis syn_module_defined=1 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(32[13:44])
    inverter_U506 \inverter_chain_543..inv  (.\notGate[542]_keep (notGate_542), 
            .\notGate[543] (notGate_543)) /* synthesis syn_module_defined=1 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(32[13:44])
    inverter_U507 \inverter_chain_542..inv  (.\notGate[541]_keep (notGate_541), 
            .\notGate[542] (notGate_542)) /* synthesis syn_module_defined=1 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(32[13:44])
    inverter_U508 \inverter_chain_541..inv  (.\notGate[540]_keep (notGate_540), 
            .\notGate[541] (notGate_541)) /* synthesis syn_module_defined=1 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(32[13:44])
    inverter_U509 \inverter_chain_540..inv  (.\notGate[539]_keep (notGate_539), 
            .\notGate[540] (notGate_540)) /* synthesis syn_module_defined=1 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(32[13:44])
    inverter_U510 \inverter_chain_53..inv  (.\notGate[52]_keep (notGate_52), 
            .\notGate[53] (notGate_53)) /* synthesis syn_module_defined=1 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(32[13:44])
    inverter_U511 \inverter_chain_539..inv  (.\notGate[538]_keep (notGate_538), 
            .\notGate[539] (notGate_539)) /* synthesis syn_module_defined=1 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(32[13:44])
    inverter_U512 \inverter_chain_538..inv  (.\notGate[537]_keep (notGate_537), 
            .\notGate[538] (notGate_538)) /* synthesis syn_module_defined=1 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(32[13:44])
    inverter_U513 \inverter_chain_537..inv  (.\notGate[536]_keep (notGate_536), 
            .\notGate[537] (notGate_537)) /* synthesis syn_module_defined=1 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(32[13:44])
    inverter_U514 \inverter_chain_536..inv  (.\notGate[535]_keep (notGate_535), 
            .\notGate[536] (notGate_536)) /* synthesis syn_module_defined=1 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(32[13:44])
    inverter_U515 \inverter_chain_535..inv  (.\notGate[534]_keep (notGate_534), 
            .\notGate[535] (notGate_535)) /* synthesis syn_module_defined=1 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(32[13:44])
    inverter_U516 \inverter_chain_534..inv  (.\notGate[533]_keep (notGate_533), 
            .\notGate[534] (notGate_534)) /* synthesis syn_module_defined=1 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(32[13:44])
    inverter_U517 \inverter_chain_533..inv  (.\notGate[532]_keep (notGate_532), 
            .\notGate[533] (notGate_533)) /* synthesis syn_module_defined=1 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(32[13:44])
    inverter_U518 \inverter_chain_532..inv  (.\notGate[531]_keep (notGate_531), 
            .\notGate[532] (notGate_532)) /* synthesis syn_module_defined=1 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(32[13:44])
    inverter_U519 \inverter_chain_531..inv  (.\notGate[530]_keep (notGate_530), 
            .\notGate[531] (notGate_531)) /* synthesis syn_module_defined=1 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(32[13:44])
    inverter_U520 \inverter_chain_530..inv  (.\notGate[529]_keep (notGate_529), 
            .\notGate[530] (notGate_530)) /* synthesis syn_module_defined=1 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(32[13:44])
    inverter_U521 \inverter_chain_52..inv  (.\notGate[51]_keep (notGate_51), 
            .\notGate[52] (notGate_52)) /* synthesis syn_module_defined=1 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(32[13:44])
    inverter_U522 \inverter_chain_529..inv  (.\notGate[528]_keep (notGate_528), 
            .\notGate[529] (notGate_529)) /* synthesis syn_module_defined=1 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(32[13:44])
    inverter_U523 \inverter_chain_528..inv  (.\notGate[527]_keep (notGate_527), 
            .\notGate[528] (notGate_528)) /* synthesis syn_module_defined=1 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(32[13:44])
    inverter_U524 \inverter_chain_527..inv  (.\notGate[526]_keep (notGate_526), 
            .\notGate[527] (notGate_527)) /* synthesis syn_module_defined=1 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(32[13:44])
    inverter_U525 \inverter_chain_526..inv  (.\notGate[525]_keep (notGate_525), 
            .\notGate[526] (notGate_526)) /* synthesis syn_module_defined=1 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(32[13:44])
    inverter_U526 \inverter_chain_525..inv  (.\notGate[524]_keep (notGate_524), 
            .\notGate[525] (notGate_525)) /* synthesis syn_module_defined=1 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(32[13:44])
    inverter_U527 \inverter_chain_524..inv  (.\notGate[523]_keep (notGate_523), 
            .\notGate[524] (notGate_524)) /* synthesis syn_module_defined=1 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(32[13:44])
    inverter_U528 \inverter_chain_523..inv  (.\notGate[522]_keep (notGate_522), 
            .\notGate[523] (notGate_523)) /* synthesis syn_module_defined=1 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(32[13:44])
    inverter_U529 \inverter_chain_522..inv  (.\notGate[521]_keep (notGate_521), 
            .\notGate[522] (notGate_522)) /* synthesis syn_module_defined=1 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(32[13:44])
    inverter_U530 \inverter_chain_521..inv  (.\notGate[520]_keep (notGate_520), 
            .\notGate[521] (notGate_521)) /* synthesis syn_module_defined=1 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(32[13:44])
    inverter_U531 \inverter_chain_520..inv  (.\notGate[519]_keep (notGate_519), 
            .\notGate[520] (notGate_520)) /* synthesis syn_module_defined=1 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(32[13:44])
    inverter_U532 \inverter_chain_51..inv  (.\notGate[50]_keep (notGate_50), 
            .\notGate[51] (notGate_51)) /* synthesis syn_module_defined=1 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(32[13:44])
    inverter_U533 \inverter_chain_519..inv  (.\notGate[518]_keep (notGate_518), 
            .\notGate[519] (notGate_519)) /* synthesis syn_module_defined=1 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(32[13:44])
    inverter_U534 \inverter_chain_518..inv  (.\notGate[517]_keep (notGate_517), 
            .\notGate[518] (notGate_518)) /* synthesis syn_module_defined=1 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(32[13:44])
    inverter_U535 \inverter_chain_517..inv  (.\notGate[516]_keep (notGate_516), 
            .\notGate[517] (notGate_517)) /* synthesis syn_module_defined=1 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(32[13:44])
    inverter_U536 \inverter_chain_516..inv  (.\notGate[515]_keep (notGate_515), 
            .\notGate[516] (notGate_516)) /* synthesis syn_module_defined=1 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(32[13:44])
    inverter_U537 \inverter_chain_515..inv  (.\notGate[514]_keep (notGate_514), 
            .\notGate[515] (notGate_515)) /* synthesis syn_module_defined=1 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(32[13:44])
    inverter_U538 \inverter_chain_514..inv  (.\notGate[513]_keep (notGate_513), 
            .\notGate[514] (notGate_514)) /* synthesis syn_module_defined=1 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(32[13:44])
    inverter_U539 \inverter_chain_513..inv  (.\notGate[512]_keep (notGate_512), 
            .\notGate[513] (notGate_513)) /* synthesis syn_module_defined=1 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(32[13:44])
    inverter_U540 \inverter_chain_512..inv  (.\notGate[511]_keep (notGate_511), 
            .\notGate[512] (notGate_512)) /* synthesis syn_module_defined=1 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(32[13:44])
    inverter_U541 \inverter_chain_511..inv  (.\notGate[510]_keep (notGate_510), 
            .\notGate[511] (notGate_511)) /* synthesis syn_module_defined=1 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(32[13:44])
    inverter_U542 \inverter_chain_510..inv  (.\notGate[509]_keep (notGate_509), 
            .\notGate[510] (notGate_510)) /* synthesis syn_module_defined=1 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(32[13:44])
    inverter_U543 \inverter_chain_50..inv  (.\notGate[49]_keep (notGate_49), 
            .\notGate[50] (notGate_50)) /* synthesis syn_module_defined=1 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(32[13:44])
    inverter_U544 \inverter_chain_509..inv  (.\notGate[508]_keep (notGate_508), 
            .\notGate[509] (notGate_509)) /* synthesis syn_module_defined=1 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(32[13:44])
    inverter_U545 \inverter_chain_508..inv  (.\notGate[507]_keep (notGate_507), 
            .\notGate[508] (notGate_508)) /* synthesis syn_module_defined=1 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(32[13:44])
    inverter_U546 \inverter_chain_507..inv  (.\notGate[506]_keep (notGate_506), 
            .\notGate[507] (notGate_507)) /* synthesis syn_module_defined=1 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(32[13:44])
    inverter_U547 \inverter_chain_506..inv  (.\notGate[505]_keep (notGate_505), 
            .\notGate[506] (notGate_506)) /* synthesis syn_module_defined=1 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(32[13:44])
    inverter_U548 \inverter_chain_505..inv  (.\notGate[504]_keep (notGate_504), 
            .\notGate[505] (notGate_505)) /* synthesis syn_module_defined=1 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(32[13:44])
    inverter_U549 \inverter_chain_504..inv  (.\notGate[503]_keep (notGate_503), 
            .\notGate[504] (notGate_504)) /* synthesis syn_module_defined=1 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(32[13:44])
    inverter_U550 \inverter_chain_503..inv  (.\notGate[502]_keep (notGate_502), 
            .\notGate[503] (notGate_503)) /* synthesis syn_module_defined=1 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(32[13:44])
    inverter_U551 \inverter_chain_502..inv  (.\notGate[501]_keep (notGate_501), 
            .\notGate[502] (notGate_502)) /* synthesis syn_module_defined=1 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(32[13:44])
    inverter_U552 \inverter_chain_501..inv  (.\notGate[500]_keep (notGate_500), 
            .\notGate[501] (notGate_501)) /* synthesis syn_module_defined=1 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(32[13:44])
    inverter_U553 \inverter_chain_500..inv  (.\notGate[499]_keep (notGate_499), 
            .\notGate[500] (notGate_500)) /* synthesis syn_module_defined=1 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(32[13:44])
    inverter_U554 \inverter_chain_4..inv  (.\notGate[3]_keep (notGate_3), 
            .\notGate[4] (notGate_4)) /* synthesis syn_module_defined=1 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(32[13:44])
    inverter_U555 \inverter_chain_49..inv  (.\notGate[48]_keep (notGate_48), 
            .\notGate[49] (notGate_49)) /* synthesis syn_module_defined=1 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(32[13:44])
    inverter_U556 \inverter_chain_499..inv  (.\notGate[498]_keep (notGate_498), 
            .\notGate[499] (notGate_499)) /* synthesis syn_module_defined=1 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(32[13:44])
    inverter_U557 \inverter_chain_498..inv  (.\notGate[497]_keep (notGate_497), 
            .\notGate[498] (notGate_498)) /* synthesis syn_module_defined=1 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(32[13:44])
    inverter_U558 \inverter_chain_497..inv  (.\notGate[496]_keep (notGate_496), 
            .\notGate[497] (notGate_497)) /* synthesis syn_module_defined=1 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(32[13:44])
    inverter_U559 \inverter_chain_496..inv  (.\notGate[495]_keep (notGate_495), 
            .\notGate[496] (notGate_496)) /* synthesis syn_module_defined=1 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(32[13:44])
    inverter_U560 \inverter_chain_495..inv  (.\notGate[494]_keep (notGate_494), 
            .\notGate[495] (notGate_495)) /* synthesis syn_module_defined=1 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(32[13:44])
    inverter_U561 \inverter_chain_494..inv  (.\notGate[493]_keep (notGate_493), 
            .\notGate[494] (notGate_494)) /* synthesis syn_module_defined=1 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(32[13:44])
    inverter_U562 \inverter_chain_493..inv  (.\notGate[492]_keep (notGate_492), 
            .\notGate[493] (notGate_493)) /* synthesis syn_module_defined=1 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(32[13:44])
    inverter_U563 \inverter_chain_492..inv  (.\notGate[491]_keep (notGate_491), 
            .\notGate[492] (notGate_492)) /* synthesis syn_module_defined=1 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(32[13:44])
    inverter_U564 \inverter_chain_491..inv  (.\notGate[490]_keep (notGate_490), 
            .\notGate[491] (notGate_491)) /* synthesis syn_module_defined=1 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(32[13:44])
    inverter_U565 \inverter_chain_490..inv  (.\notGate[489]_keep (notGate_489), 
            .\notGate[490] (notGate_490)) /* synthesis syn_module_defined=1 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(32[13:44])
    inverter_U566 \inverter_chain_48..inv  (.\notGate[47]_keep (notGate_47), 
            .\notGate[48] (notGate_48)) /* synthesis syn_module_defined=1 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(32[13:44])
    inverter_U567 \inverter_chain_489..inv  (.\notGate[488]_keep (notGate_488), 
            .\notGate[489] (notGate_489)) /* synthesis syn_module_defined=1 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(32[13:44])
    inverter_U568 \inverter_chain_488..inv  (.\notGate[487]_keep (notGate_487), 
            .\notGate[488] (notGate_488)) /* synthesis syn_module_defined=1 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(32[13:44])
    inverter_U569 \inverter_chain_487..inv  (.\notGate[486]_keep (notGate_486), 
            .\notGate[487] (notGate_487)) /* synthesis syn_module_defined=1 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(32[13:44])
    inverter_U570 \inverter_chain_486..inv  (.\notGate[485]_keep (notGate_485), 
            .\notGate[486] (notGate_486)) /* synthesis syn_module_defined=1 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(32[13:44])
    inverter_U571 \inverter_chain_485..inv  (.\notGate[484]_keep (notGate_484), 
            .\notGate[485] (notGate_485)) /* synthesis syn_module_defined=1 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(32[13:44])
    inverter_U572 \inverter_chain_484..inv  (.\notGate[483]_keep (notGate_483), 
            .\notGate[484] (notGate_484)) /* synthesis syn_module_defined=1 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(32[13:44])
    inverter_U573 \inverter_chain_483..inv  (.\notGate[482]_keep (notGate_482), 
            .\notGate[483] (notGate_483)) /* synthesis syn_module_defined=1 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(32[13:44])
    inverter_U574 \inverter_chain_482..inv  (.\notGate[481]_keep (notGate_481), 
            .\notGate[482] (notGate_482)) /* synthesis syn_module_defined=1 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(32[13:44])
    inverter_U575 \inverter_chain_481..inv  (.\notGate[480]_keep (notGate_480), 
            .\notGate[481] (notGate_481)) /* synthesis syn_module_defined=1 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(32[13:44])
    inverter_U576 \inverter_chain_480..inv  (.\notGate[479]_keep (notGate_479), 
            .\notGate[480] (notGate_480)) /* synthesis syn_module_defined=1 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(32[13:44])
    inverter_U577 \inverter_chain_47..inv  (.\notGate[46]_keep (notGate_46), 
            .\notGate[47] (notGate_47)) /* synthesis syn_module_defined=1 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(32[13:44])
    inverter_U578 \inverter_chain_479..inv  (.\notGate[478]_keep (notGate_478), 
            .\notGate[479] (notGate_479)) /* synthesis syn_module_defined=1 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(32[13:44])
    inverter_U579 \inverter_chain_478..inv  (.\notGate[477]_keep (notGate_477), 
            .\notGate[478] (notGate_478)) /* synthesis syn_module_defined=1 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(32[13:44])
    inverter_U580 \inverter_chain_477..inv  (.\notGate[476]_keep (notGate_476), 
            .\notGate[477] (notGate_477)) /* synthesis syn_module_defined=1 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(32[13:44])
    inverter_U581 \inverter_chain_476..inv  (.\notGate[475]_keep (notGate_475), 
            .\notGate[476] (notGate_476)) /* synthesis syn_module_defined=1 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(32[13:44])
    inverter_U582 \inverter_chain_475..inv  (.\notGate[474]_keep (notGate_474), 
            .\notGate[475] (notGate_475)) /* synthesis syn_module_defined=1 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(32[13:44])
    inverter_U583 \inverter_chain_474..inv  (.\notGate[473]_keep (notGate_473), 
            .\notGate[474] (notGate_474)) /* synthesis syn_module_defined=1 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(32[13:44])
    inverter_U584 \inverter_chain_473..inv  (.\notGate[472]_keep (notGate_472), 
            .\notGate[473] (notGate_473)) /* synthesis syn_module_defined=1 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(32[13:44])
    inverter_U585 \inverter_chain_472..inv  (.\notGate[471]_keep (notGate_471), 
            .\notGate[472] (notGate_472)) /* synthesis syn_module_defined=1 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(32[13:44])
    inverter_U586 \inverter_chain_471..inv  (.\notGate[470]_keep (notGate_470), 
            .\notGate[471] (notGate_471)) /* synthesis syn_module_defined=1 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(32[13:44])
    inverter_U587 \inverter_chain_470..inv  (.\notGate[469]_keep (notGate_469), 
            .\notGate[470] (notGate_470)) /* synthesis syn_module_defined=1 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(32[13:44])
    inverter_U588 \inverter_chain_46..inv  (.\notGate[45]_keep (notGate_45), 
            .\notGate[46] (notGate_46)) /* synthesis syn_module_defined=1 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(32[13:44])
    inverter_U589 \inverter_chain_469..inv  (.\notGate[468]_keep (notGate_468), 
            .\notGate[469] (notGate_469)) /* synthesis syn_module_defined=1 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(32[13:44])
    inverter_U590 \inverter_chain_468..inv  (.\notGate[467]_keep (notGate_467), 
            .\notGate[468] (notGate_468)) /* synthesis syn_module_defined=1 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(32[13:44])
    inverter_U591 \inverter_chain_467..inv  (.\notGate[466]_keep (notGate_466), 
            .\notGate[467] (notGate_467)) /* synthesis syn_module_defined=1 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(32[13:44])
    inverter_U592 \inverter_chain_466..inv  (.\notGate[465]_keep (notGate_465), 
            .\notGate[466] (notGate_466)) /* synthesis syn_module_defined=1 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(32[13:44])
    inverter_U593 \inverter_chain_465..inv  (.\notGate[464]_keep (notGate_464), 
            .\notGate[465] (notGate_465)) /* synthesis syn_module_defined=1 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(32[13:44])
    inverter_U594 \inverter_chain_464..inv  (.\notGate[463]_keep (notGate_463), 
            .\notGate[464] (notGate_464)) /* synthesis syn_module_defined=1 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(32[13:44])
    inverter_U595 \inverter_chain_463..inv  (.\notGate[462]_keep (notGate_462), 
            .\notGate[463] (notGate_463)) /* synthesis syn_module_defined=1 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(32[13:44])
    inverter_U596 \inverter_chain_462..inv  (.\notGate[461]_keep (notGate_461), 
            .\notGate[462] (notGate_462)) /* synthesis syn_module_defined=1 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(32[13:44])
    inverter_U597 \inverter_chain_461..inv  (.\notGate[460]_keep (notGate_460), 
            .\notGate[461] (notGate_461)) /* synthesis syn_module_defined=1 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(32[13:44])
    inverter_U598 \inverter_chain_460..inv  (.\notGate[459]_keep (notGate_459), 
            .\notGate[460] (notGate_460)) /* synthesis syn_module_defined=1 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(32[13:44])
    inverter_U599 \inverter_chain_45..inv  (.\notGate[44]_keep (notGate_44), 
            .\notGate[45] (notGate_45)) /* synthesis syn_module_defined=1 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(32[13:44])
    inverter_U600 \inverter_chain_459..inv  (.\notGate[458]_keep (notGate_458), 
            .\notGate[459] (notGate_459)) /* synthesis syn_module_defined=1 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(32[13:44])
    inverter_U601 \inverter_chain_458..inv  (.\notGate[457]_keep (notGate_457), 
            .\notGate[458] (notGate_458)) /* synthesis syn_module_defined=1 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(32[13:44])
    inverter_U602 \inverter_chain_457..inv  (.\notGate[456]_keep (notGate_456), 
            .\notGate[457] (notGate_457)) /* synthesis syn_module_defined=1 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(32[13:44])
    inverter_U603 \inverter_chain_456..inv  (.\notGate[455]_keep (notGate_455), 
            .\notGate[456] (notGate_456)) /* synthesis syn_module_defined=1 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(32[13:44])
    inverter_U604 \inverter_chain_455..inv  (.\notGate[454]_keep (notGate_454), 
            .\notGate[455] (notGate_455)) /* synthesis syn_module_defined=1 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(32[13:44])
    inverter_U605 \inverter_chain_454..inv  (.\notGate[453]_keep (notGate_453), 
            .\notGate[454] (notGate_454)) /* synthesis syn_module_defined=1 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(32[13:44])
    inverter_U606 \inverter_chain_453..inv  (.\notGate[452]_keep (notGate_452), 
            .\notGate[453] (notGate_453)) /* synthesis syn_module_defined=1 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(32[13:44])
    inverter_U607 \inverter_chain_452..inv  (.\notGate[451]_keep (notGate_451), 
            .\notGate[452] (notGate_452)) /* synthesis syn_module_defined=1 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(32[13:44])
    inverter_U608 \inverter_chain_451..inv  (.\notGate[450]_keep (notGate_450), 
            .\notGate[451] (notGate_451)) /* synthesis syn_module_defined=1 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(32[13:44])
    inverter_U609 \inverter_chain_450..inv  (.\notGate[449]_keep (notGate_449), 
            .\notGate[450] (notGate_450)) /* synthesis syn_module_defined=1 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(32[13:44])
    inverter_U610 \inverter_chain_44..inv  (.\notGate[43]_keep (notGate_43), 
            .\notGate[44] (notGate_44)) /* synthesis syn_module_defined=1 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(32[13:44])
    inverter_U611 \inverter_chain_449..inv  (.\notGate[448]_keep (notGate_448), 
            .\notGate[449] (notGate_449)) /* synthesis syn_module_defined=1 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(32[13:44])
    inverter_U612 \inverter_chain_448..inv  (.\notGate[447]_keep (notGate_447), 
            .\notGate[448] (notGate_448)) /* synthesis syn_module_defined=1 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(32[13:44])
    inverter_U613 \inverter_chain_447..inv  (.\notGate[446]_keep (notGate_446), 
            .\notGate[447] (notGate_447)) /* synthesis syn_module_defined=1 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(32[13:44])
    inverter_U614 \inverter_chain_446..inv  (.\notGate[445]_keep (notGate_445), 
            .\notGate[446] (notGate_446)) /* synthesis syn_module_defined=1 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(32[13:44])
    inverter_U615 \inverter_chain_445..inv  (.\notGate[444]_keep (notGate_444), 
            .\notGate[445] (notGate_445)) /* synthesis syn_module_defined=1 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(32[13:44])
    inverter_U616 \inverter_chain_444..inv  (.\notGate[443]_keep (notGate_443), 
            .\notGate[444] (notGate_444)) /* synthesis syn_module_defined=1 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(32[13:44])
    inverter_U617 \inverter_chain_443..inv  (.\notGate[442]_keep (notGate_442), 
            .\notGate[443] (notGate_443)) /* synthesis syn_module_defined=1 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(32[13:44])
    inverter_U618 \inverter_chain_442..inv  (.\notGate[441]_keep (notGate_441), 
            .\notGate[442] (notGate_442)) /* synthesis syn_module_defined=1 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(32[13:44])
    inverter_U619 \inverter_chain_441..inv  (.\notGate[440]_keep (notGate_440), 
            .\notGate[441] (notGate_441)) /* synthesis syn_module_defined=1 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(32[13:44])
    inverter_U620 \inverter_chain_440..inv  (.\notGate[439]_keep (notGate_439), 
            .\notGate[440] (notGate_440)) /* synthesis syn_module_defined=1 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(32[13:44])
    inverter_U621 \inverter_chain_43..inv  (.\notGate[42]_keep (notGate_42), 
            .\notGate[43] (notGate_43)) /* synthesis syn_module_defined=1 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(32[13:44])
    inverter_U622 \inverter_chain_439..inv  (.\notGate[438]_keep (notGate_438), 
            .\notGate[439] (notGate_439)) /* synthesis syn_module_defined=1 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(32[13:44])
    inverter_U623 \inverter_chain_438..inv  (.\notGate[437]_keep (notGate_437), 
            .\notGate[438] (notGate_438)) /* synthesis syn_module_defined=1 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(32[13:44])
    inverter_U624 \inverter_chain_437..inv  (.\notGate[436]_keep (notGate_436), 
            .\notGate[437] (notGate_437)) /* synthesis syn_module_defined=1 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(32[13:44])
    inverter_U625 \inverter_chain_436..inv  (.\notGate[435]_keep (notGate_435), 
            .\notGate[436] (notGate_436)) /* synthesis syn_module_defined=1 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(32[13:44])
    inverter_U626 \inverter_chain_435..inv  (.\notGate[434]_keep (notGate_434), 
            .\notGate[435] (notGate_435)) /* synthesis syn_module_defined=1 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(32[13:44])
    inverter_U627 \inverter_chain_434..inv  (.\notGate[433]_keep (notGate_433), 
            .\notGate[434] (notGate_434)) /* synthesis syn_module_defined=1 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(32[13:44])
    inverter_U628 \inverter_chain_433..inv  (.\notGate[432]_keep (notGate_432), 
            .\notGate[433] (notGate_433)) /* synthesis syn_module_defined=1 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(32[13:44])
    inverter_U629 \inverter_chain_432..inv  (.\notGate[431]_keep (notGate_431), 
            .\notGate[432] (notGate_432)) /* synthesis syn_module_defined=1 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(32[13:44])
    inverter_U630 \inverter_chain_431..inv  (.\notGate[430]_keep (notGate_430), 
            .\notGate[431] (notGate_431)) /* synthesis syn_module_defined=1 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(32[13:44])
    inverter_U631 \inverter_chain_430..inv  (.\notGate[429]_keep (notGate_429), 
            .\notGate[430] (notGate_430)) /* synthesis syn_module_defined=1 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(32[13:44])
    inverter_U632 \inverter_chain_42..inv  (.\notGate[41]_keep (notGate_41), 
            .\notGate[42] (notGate_42)) /* synthesis syn_module_defined=1 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(32[13:44])
    inverter_U633 \inverter_chain_429..inv  (.\notGate[428]_keep (notGate_428), 
            .\notGate[429] (notGate_429)) /* synthesis syn_module_defined=1 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(32[13:44])
    inverter_U634 \inverter_chain_428..inv  (.\notGate[427]_keep (notGate_427), 
            .\notGate[428] (notGate_428)) /* synthesis syn_module_defined=1 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(32[13:44])
    inverter_U635 \inverter_chain_427..inv  (.\notGate[426]_keep (notGate_426), 
            .\notGate[427] (notGate_427)) /* synthesis syn_module_defined=1 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(32[13:44])
    inverter_U636 \inverter_chain_426..inv  (.\notGate[425]_keep (notGate_425), 
            .\notGate[426] (notGate_426)) /* synthesis syn_module_defined=1 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(32[13:44])
    inverter_U637 \inverter_chain_425..inv  (.\notGate[424]_keep (notGate_424), 
            .\notGate[425] (notGate_425)) /* synthesis syn_module_defined=1 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(32[13:44])
    inverter_U638 \inverter_chain_424..inv  (.\notGate[423]_keep (notGate_423), 
            .\notGate[424] (notGate_424)) /* synthesis syn_module_defined=1 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(32[13:44])
    inverter_U639 \inverter_chain_423..inv  (.\notGate[422]_keep (notGate_422), 
            .\notGate[423] (notGate_423)) /* synthesis syn_module_defined=1 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(32[13:44])
    inverter_U640 \inverter_chain_422..inv  (.\notGate[421]_keep (notGate_421), 
            .\notGate[422] (notGate_422)) /* synthesis syn_module_defined=1 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(32[13:44])
    inverter_U641 \inverter_chain_421..inv  (.\notGate[420]_keep (notGate_420), 
            .\notGate[421] (notGate_421)) /* synthesis syn_module_defined=1 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(32[13:44])
    inverter_U642 \inverter_chain_420..inv  (.\notGate[419]_keep (notGate_419), 
            .\notGate[420] (notGate_420)) /* synthesis syn_module_defined=1 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(32[13:44])
    inverter_U643 \inverter_chain_41..inv  (.\notGate[40]_keep (notGate_40), 
            .\notGate[41] (notGate_41)) /* synthesis syn_module_defined=1 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(32[13:44])
    inverter_U644 \inverter_chain_419..inv  (.\notGate[418]_keep (notGate_418), 
            .\notGate[419] (notGate_419)) /* synthesis syn_module_defined=1 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(32[13:44])
    inverter_U645 \inverter_chain_418..inv  (.\notGate[417]_keep (notGate_417), 
            .\notGate[418] (notGate_418)) /* synthesis syn_module_defined=1 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(32[13:44])
    inverter_U646 \inverter_chain_417..inv  (.\notGate[416]_keep (notGate_416), 
            .\notGate[417] (notGate_417)) /* synthesis syn_module_defined=1 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(32[13:44])
    inverter_U647 \inverter_chain_416..inv  (.\notGate[415]_keep (notGate_415), 
            .\notGate[416] (notGate_416)) /* synthesis syn_module_defined=1 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(32[13:44])
    inverter_U648 \inverter_chain_415..inv  (.\notGate[414]_keep (notGate_414), 
            .\notGate[415] (notGate_415)) /* synthesis syn_module_defined=1 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(32[13:44])
    inverter_U649 \inverter_chain_414..inv  (.\notGate[413]_keep (notGate_413), 
            .\notGate[414] (notGate_414)) /* synthesis syn_module_defined=1 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(32[13:44])
    inverter_U650 \inverter_chain_413..inv  (.\notGate[412]_keep (notGate_412), 
            .\notGate[413] (notGate_413)) /* synthesis syn_module_defined=1 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(32[13:44])
    inverter_U651 \inverter_chain_412..inv  (.\notGate[411]_keep (notGate_411), 
            .\notGate[412] (notGate_412)) /* synthesis syn_module_defined=1 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(32[13:44])
    inverter_U652 \inverter_chain_411..inv  (.\notGate[410]_keep (notGate_410), 
            .\notGate[411] (notGate_411)) /* synthesis syn_module_defined=1 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(32[13:44])
    inverter_U653 \inverter_chain_410..inv  (.\notGate[409]_keep (notGate_409), 
            .\notGate[410] (notGate_410)) /* synthesis syn_module_defined=1 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(32[13:44])
    inverter_U654 \inverter_chain_40..inv  (.\notGate[39]_keep (notGate_39), 
            .\notGate[40] (notGate_40)) /* synthesis syn_module_defined=1 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(32[13:44])
    inverter_U655 \inverter_chain_409..inv  (.\notGate[408]_keep (notGate_408), 
            .\notGate[409] (notGate_409)) /* synthesis syn_module_defined=1 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(32[13:44])
    inverter_U656 \inverter_chain_408..inv  (.\notGate[407]_keep (notGate_407), 
            .\notGate[408] (notGate_408)) /* synthesis syn_module_defined=1 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(32[13:44])
    inverter_U657 \inverter_chain_407..inv  (.\notGate[406]_keep (notGate_406), 
            .\notGate[407] (notGate_407)) /* synthesis syn_module_defined=1 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(32[13:44])
    inverter_U658 \inverter_chain_406..inv  (.\notGate[405]_keep (notGate_405), 
            .\notGate[406] (notGate_406)) /* synthesis syn_module_defined=1 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(32[13:44])
    inverter_U659 \inverter_chain_405..inv  (.\notGate[404]_keep (notGate_404), 
            .\notGate[405] (notGate_405)) /* synthesis syn_module_defined=1 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(32[13:44])
    inverter_U660 \inverter_chain_404..inv  (.\notGate[403]_keep (notGate_403), 
            .\notGate[404] (notGate_404)) /* synthesis syn_module_defined=1 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(32[13:44])
    inverter_U661 \inverter_chain_403..inv  (.\notGate[402]_keep (notGate_402), 
            .\notGate[403] (notGate_403)) /* synthesis syn_module_defined=1 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(32[13:44])
    inverter_U662 \inverter_chain_402..inv  (.\notGate[401]_keep (notGate_401), 
            .\notGate[402] (notGate_402)) /* synthesis syn_module_defined=1 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(32[13:44])
    inverter_U663 \inverter_chain_401..inv  (.\notGate[400]_keep (notGate_400), 
            .\notGate[401] (notGate_401)) /* synthesis syn_module_defined=1 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(32[13:44])
    inverter_U664 \inverter_chain_400..inv  (.\notGate[399]_keep (notGate_399), 
            .\notGate[400] (notGate_400)) /* synthesis syn_module_defined=1 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(32[13:44])
    inverter_U665 \inverter_chain_3..inv  (.\notGate[2]_keep (notGate_2), 
            .\notGate[3] (notGate_3)) /* synthesis syn_module_defined=1 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(32[13:44])
    inverter_U666 \inverter_chain_39..inv  (.\notGate[38]_keep (notGate_38), 
            .\notGate[39] (notGate_39)) /* synthesis syn_module_defined=1 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(32[13:44])
    inverter_U667 \inverter_chain_399..inv  (.\notGate[398]_keep (notGate_398), 
            .\notGate[399] (notGate_399)) /* synthesis syn_module_defined=1 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(32[13:44])
    inverter_U668 \inverter_chain_398..inv  (.\notGate[397]_keep (notGate_397), 
            .\notGate[398] (notGate_398)) /* synthesis syn_module_defined=1 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(32[13:44])
    inverter_U669 \inverter_chain_397..inv  (.\notGate[396]_keep (notGate_396), 
            .\notGate[397] (notGate_397)) /* synthesis syn_module_defined=1 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(32[13:44])
    inverter_U670 \inverter_chain_396..inv  (.\notGate[395]_keep (notGate_395), 
            .\notGate[396] (notGate_396)) /* synthesis syn_module_defined=1 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(32[13:44])
    inverter_U671 \inverter_chain_395..inv  (.\notGate[394]_keep (notGate_394), 
            .\notGate[395] (notGate_395)) /* synthesis syn_module_defined=1 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(32[13:44])
    inverter_U672 \inverter_chain_394..inv  (.\notGate[393]_keep (notGate_393), 
            .\notGate[394] (notGate_394)) /* synthesis syn_module_defined=1 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(32[13:44])
    inverter_U673 \inverter_chain_393..inv  (.\notGate[392]_keep (notGate_392), 
            .\notGate[393] (notGate_393)) /* synthesis syn_module_defined=1 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(32[13:44])
    inverter_U674 \inverter_chain_392..inv  (.\notGate[391]_keep (notGate_391), 
            .\notGate[392] (notGate_392)) /* synthesis syn_module_defined=1 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(32[13:44])
    inverter_U675 \inverter_chain_391..inv  (.\notGate[390]_keep (notGate_390), 
            .\notGate[391] (notGate_391)) /* synthesis syn_module_defined=1 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(32[13:44])
    inverter_U676 \inverter_chain_390..inv  (.\notGate[389]_keep (notGate_389), 
            .\notGate[390] (notGate_390)) /* synthesis syn_module_defined=1 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(32[13:44])
    inverter_U677 \inverter_chain_38..inv  (.\notGate[37]_keep (notGate_37), 
            .\notGate[38] (notGate_38)) /* synthesis syn_module_defined=1 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(32[13:44])
    inverter_U678 \inverter_chain_389..inv  (.\notGate[388]_keep (notGate_388), 
            .\notGate[389] (notGate_389)) /* synthesis syn_module_defined=1 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(32[13:44])
    inverter_U679 \inverter_chain_388..inv  (.\notGate[387]_keep (notGate_387), 
            .\notGate[388] (notGate_388)) /* synthesis syn_module_defined=1 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(32[13:44])
    inverter_U680 \inverter_chain_387..inv  (.\notGate[386]_keep (notGate_386), 
            .\notGate[387] (notGate_387)) /* synthesis syn_module_defined=1 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(32[13:44])
    inverter_U681 \inverter_chain_386..inv  (.\notGate[385]_keep (notGate_385), 
            .\notGate[386] (notGate_386)) /* synthesis syn_module_defined=1 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(32[13:44])
    inverter_U682 \inverter_chain_385..inv  (.\notGate[384]_keep (notGate_384), 
            .\notGate[385] (notGate_385)) /* synthesis syn_module_defined=1 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(32[13:44])
    inverter_U683 \inverter_chain_384..inv  (.\notGate[383]_keep (notGate_383), 
            .\notGate[384] (notGate_384)) /* synthesis syn_module_defined=1 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(32[13:44])
    inverter_U684 \inverter_chain_383..inv  (.\notGate[382]_keep (notGate_382), 
            .\notGate[383] (notGate_383)) /* synthesis syn_module_defined=1 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(32[13:44])
    inverter_U685 \inverter_chain_382..inv  (.\notGate[381]_keep (notGate_381), 
            .\notGate[382] (notGate_382)) /* synthesis syn_module_defined=1 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(32[13:44])
    inverter_U686 \inverter_chain_381..inv  (.\notGate[380]_keep (notGate_380), 
            .\notGate[381] (notGate_381)) /* synthesis syn_module_defined=1 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(32[13:44])
    inverter_U687 \inverter_chain_380..inv  (.\notGate[379]_keep (notGate_379), 
            .\notGate[380] (notGate_380)) /* synthesis syn_module_defined=1 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(32[13:44])
    inverter_U688 \inverter_chain_37..inv  (.\notGate[36]_keep (notGate_36), 
            .\notGate[37] (notGate_37)) /* synthesis syn_module_defined=1 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(32[13:44])
    inverter_U689 \inverter_chain_379..inv  (.\notGate[378]_keep (notGate_378), 
            .\notGate[379] (notGate_379)) /* synthesis syn_module_defined=1 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(32[13:44])
    inverter_U690 \inverter_chain_378..inv  (.\notGate[377]_keep (notGate_377), 
            .\notGate[378] (notGate_378)) /* synthesis syn_module_defined=1 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(32[13:44])
    inverter_U691 \inverter_chain_377..inv  (.\notGate[376]_keep (notGate_376), 
            .\notGate[377] (notGate_377)) /* synthesis syn_module_defined=1 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(32[13:44])
    inverter_U692 \inverter_chain_376..inv  (.\notGate[375]_keep (notGate_375), 
            .\notGate[376] (notGate_376)) /* synthesis syn_module_defined=1 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(32[13:44])
    inverter_U693 \inverter_chain_375..inv  (.\notGate[374]_keep (notGate_374), 
            .\notGate[375] (notGate_375)) /* synthesis syn_module_defined=1 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(32[13:44])
    inverter_U694 \inverter_chain_374..inv  (.\notGate[373]_keep (notGate_373), 
            .\notGate[374] (notGate_374)) /* synthesis syn_module_defined=1 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(32[13:44])
    inverter_U695 \inverter_chain_373..inv  (.\notGate[372]_keep (notGate_372), 
            .\notGate[373] (notGate_373)) /* synthesis syn_module_defined=1 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(32[13:44])
    inverter_U696 \inverter_chain_372..inv  (.\notGate[371]_keep (notGate_371), 
            .\notGate[372] (notGate_372)) /* synthesis syn_module_defined=1 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(32[13:44])
    inverter_U697 \inverter_chain_371..inv  (.\notGate[370]_keep (notGate_370), 
            .\notGate[371] (notGate_371)) /* synthesis syn_module_defined=1 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(32[13:44])
    inverter_U698 \inverter_chain_370..inv  (.\notGate[369]_keep (notGate_369), 
            .\notGate[370] (notGate_370)) /* synthesis syn_module_defined=1 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(32[13:44])
    inverter_U699 \inverter_chain_36..inv  (.\notGate[35]_keep (notGate_35), 
            .\notGate[36] (notGate_36)) /* synthesis syn_module_defined=1 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(32[13:44])
    inverter_U700 \inverter_chain_369..inv  (.\notGate[368]_keep (notGate_368), 
            .\notGate[369] (notGate_369)) /* synthesis syn_module_defined=1 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(32[13:44])
    inverter_U701 \inverter_chain_368..inv  (.\notGate[367]_keep (notGate_367), 
            .\notGate[368] (notGate_368)) /* synthesis syn_module_defined=1 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(32[13:44])
    inverter_U702 \inverter_chain_367..inv  (.\notGate[366]_keep (notGate_366), 
            .\notGate[367] (notGate_367)) /* synthesis syn_module_defined=1 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(32[13:44])
    inverter_U703 \inverter_chain_366..inv  (.\notGate[365]_keep (notGate_365), 
            .\notGate[366] (notGate_366)) /* synthesis syn_module_defined=1 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(32[13:44])
    inverter_U704 \inverter_chain_365..inv  (.\notGate[364]_keep (notGate_364), 
            .\notGate[365] (notGate_365)) /* synthesis syn_module_defined=1 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(32[13:44])
    inverter_U705 \inverter_chain_364..inv  (.\notGate[363]_keep (notGate_363), 
            .\notGate[364] (notGate_364)) /* synthesis syn_module_defined=1 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(32[13:44])
    inverter_U706 \inverter_chain_363..inv  (.\notGate[362]_keep (notGate_362), 
            .\notGate[363] (notGate_363)) /* synthesis syn_module_defined=1 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(32[13:44])
    inverter_U707 \inverter_chain_362..inv  (.\notGate[361]_keep (notGate_361), 
            .\notGate[362] (notGate_362)) /* synthesis syn_module_defined=1 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(32[13:44])
    inverter_U708 \inverter_chain_361..inv  (.\notGate[360]_keep (notGate_360), 
            .\notGate[361] (notGate_361)) /* synthesis syn_module_defined=1 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(32[13:44])
    inverter_U709 \inverter_chain_360..inv  (.\notGate[359]_keep (notGate_359), 
            .\notGate[360] (notGate_360)) /* synthesis syn_module_defined=1 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(32[13:44])
    inverter_U710 \inverter_chain_35..inv  (.\notGate[34]_keep (notGate_34), 
            .\notGate[35] (notGate_35)) /* synthesis syn_module_defined=1 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(32[13:44])
    inverter_U711 \inverter_chain_359..inv  (.\notGate[358]_keep (notGate_358), 
            .\notGate[359] (notGate_359)) /* synthesis syn_module_defined=1 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(32[13:44])
    inverter_U712 \inverter_chain_358..inv  (.\notGate[357]_keep (notGate_357), 
            .\notGate[358] (notGate_358)) /* synthesis syn_module_defined=1 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(32[13:44])
    inverter_U713 \inverter_chain_357..inv  (.\notGate[356]_keep (notGate_356), 
            .\notGate[357] (notGate_357)) /* synthesis syn_module_defined=1 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(32[13:44])
    inverter_U714 \inverter_chain_356..inv  (.\notGate[355]_keep (notGate_355), 
            .\notGate[356] (notGate_356)) /* synthesis syn_module_defined=1 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(32[13:44])
    inverter_U715 \inverter_chain_355..inv  (.\notGate[354]_keep (notGate_354), 
            .\notGate[355] (notGate_355)) /* synthesis syn_module_defined=1 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(32[13:44])
    inverter_U716 \inverter_chain_354..inv  (.\notGate[353]_keep (notGate_353), 
            .\notGate[354] (notGate_354)) /* synthesis syn_module_defined=1 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(32[13:44])
    inverter_U717 \inverter_chain_353..inv  (.\notGate[352]_keep (notGate_352), 
            .\notGate[353] (notGate_353)) /* synthesis syn_module_defined=1 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(32[13:44])
    inverter_U718 \inverter_chain_352..inv  (.\notGate[351]_keep (notGate_351), 
            .\notGate[352] (notGate_352)) /* synthesis syn_module_defined=1 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(32[13:44])
    inverter_U719 \inverter_chain_351..inv  (.\notGate[350]_keep (notGate_350), 
            .\notGate[351] (notGate_351)) /* synthesis syn_module_defined=1 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(32[13:44])
    inverter_U720 \inverter_chain_350..inv  (.\notGate[349]_keep (notGate_349), 
            .\notGate[350] (notGate_350)) /* synthesis syn_module_defined=1 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(32[13:44])
    inverter_U721 \inverter_chain_34..inv  (.\notGate[33]_keep (notGate_33), 
            .\notGate[34] (notGate_34)) /* synthesis syn_module_defined=1 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(32[13:44])
    inverter_U722 \inverter_chain_349..inv  (.\notGate[348]_keep (notGate_348), 
            .\notGate[349] (notGate_349)) /* synthesis syn_module_defined=1 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(32[13:44])
    inverter_U723 \inverter_chain_348..inv  (.\notGate[347]_keep (notGate_347), 
            .\notGate[348] (notGate_348)) /* synthesis syn_module_defined=1 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(32[13:44])
    inverter_U724 \inverter_chain_347..inv  (.\notGate[346]_keep (notGate_346), 
            .\notGate[347] (notGate_347)) /* synthesis syn_module_defined=1 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(32[13:44])
    inverter_U725 \inverter_chain_346..inv  (.\notGate[345]_keep (notGate_345), 
            .\notGate[346] (notGate_346)) /* synthesis syn_module_defined=1 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(32[13:44])
    inverter_U726 \inverter_chain_345..inv  (.\notGate[344]_keep (notGate_344), 
            .\notGate[345] (notGate_345)) /* synthesis syn_module_defined=1 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(32[13:44])
    inverter_U727 \inverter_chain_344..inv  (.\notGate[343]_keep (notGate_343), 
            .\notGate[344] (notGate_344)) /* synthesis syn_module_defined=1 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(32[13:44])
    inverter_U728 \inverter_chain_343..inv  (.\notGate[342]_keep (notGate_342), 
            .\notGate[343] (notGate_343)) /* synthesis syn_module_defined=1 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(32[13:44])
    inverter_U729 \inverter_chain_342..inv  (.\notGate[341]_keep (notGate_341), 
            .\notGate[342] (notGate_342)) /* synthesis syn_module_defined=1 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(32[13:44])
    inverter_U730 \inverter_chain_341..inv  (.\notGate[340]_keep (notGate_340), 
            .\notGate[341] (notGate_341)) /* synthesis syn_module_defined=1 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(32[13:44])
    inverter_U731 \inverter_chain_340..inv  (.\notGate[339]_keep (notGate_339), 
            .\notGate[340] (notGate_340)) /* synthesis syn_module_defined=1 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(32[13:44])
    inverter_U732 \inverter_chain_33..inv  (.\notGate[32]_keep (notGate_32), 
            .\notGate[33] (notGate_33)) /* synthesis syn_module_defined=1 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(32[13:44])
    inverter_U733 \inverter_chain_339..inv  (.\notGate[338]_keep (notGate_338), 
            .\notGate[339] (notGate_339)) /* synthesis syn_module_defined=1 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(32[13:44])
    inverter_U734 \inverter_chain_338..inv  (.\notGate[337]_keep (notGate_337), 
            .\notGate[338] (notGate_338)) /* synthesis syn_module_defined=1 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(32[13:44])
    inverter_U735 \inverter_chain_337..inv  (.\notGate[336]_keep (notGate_336), 
            .\notGate[337] (notGate_337)) /* synthesis syn_module_defined=1 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(32[13:44])
    inverter_U736 \inverter_chain_336..inv  (.\notGate[335]_keep (notGate_335), 
            .\notGate[336] (notGate_336)) /* synthesis syn_module_defined=1 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(32[13:44])
    inverter_U737 \inverter_chain_335..inv  (.\notGate[334]_keep (notGate_334), 
            .\notGate[335] (notGate_335)) /* synthesis syn_module_defined=1 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(32[13:44])
    inverter_U738 \inverter_chain_334..inv  (.\notGate[333]_keep (notGate_333), 
            .\notGate[334] (notGate_334)) /* synthesis syn_module_defined=1 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(32[13:44])
    inverter_U739 \inverter_chain_333..inv  (.\notGate[332]_keep (notGate_332), 
            .\notGate[333] (notGate_333)) /* synthesis syn_module_defined=1 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(32[13:44])
    inverter_U740 \inverter_chain_332..inv  (.\notGate[331]_keep (notGate_331), 
            .\notGate[332] (notGate_332)) /* synthesis syn_module_defined=1 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(32[13:44])
    inverter_U741 \inverter_chain_331..inv  (.\notGate[330]_keep (notGate_330), 
            .\notGate[331] (notGate_331)) /* synthesis syn_module_defined=1 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(32[13:44])
    inverter_U742 \inverter_chain_330..inv  (.\notGate[329]_keep (notGate_329), 
            .\notGate[330] (notGate_330)) /* synthesis syn_module_defined=1 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(32[13:44])
    inverter_U743 \inverter_chain_32..inv  (.\notGate[31]_keep (notGate_31), 
            .\notGate[32] (notGate_32)) /* synthesis syn_module_defined=1 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(32[13:44])
    inverter_U744 \inverter_chain_329..inv  (.\notGate[328]_keep (notGate_328), 
            .\notGate[329] (notGate_329)) /* synthesis syn_module_defined=1 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(32[13:44])
    inverter_U745 \inverter_chain_328..inv  (.\notGate[327]_keep (notGate_327), 
            .\notGate[328] (notGate_328)) /* synthesis syn_module_defined=1 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(32[13:44])
    inverter_U746 \inverter_chain_327..inv  (.\notGate[326]_keep (notGate_326), 
            .\notGate[327] (notGate_327)) /* synthesis syn_module_defined=1 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(32[13:44])
    inverter_U747 \inverter_chain_326..inv  (.\notGate[325]_keep (notGate_325), 
            .\notGate[326] (notGate_326)) /* synthesis syn_module_defined=1 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(32[13:44])
    inverter_U748 \inverter_chain_325..inv  (.\notGate[324]_keep (notGate_324), 
            .\notGate[325] (notGate_325)) /* synthesis syn_module_defined=1 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(32[13:44])
    inverter_U749 \inverter_chain_324..inv  (.\notGate[323]_keep (notGate_323), 
            .\notGate[324] (notGate_324)) /* synthesis syn_module_defined=1 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(32[13:44])
    inverter_U750 \inverter_chain_323..inv  (.\notGate[322]_keep (notGate_322), 
            .\notGate[323] (notGate_323)) /* synthesis syn_module_defined=1 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(32[13:44])
    inverter_U751 \inverter_chain_322..inv  (.\notGate[321]_keep (notGate_321), 
            .\notGate[322] (notGate_322)) /* synthesis syn_module_defined=1 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(32[13:44])
    inverter_U752 \inverter_chain_321..inv  (.\notGate[320]_keep (notGate_320), 
            .\notGate[321] (notGate_321)) /* synthesis syn_module_defined=1 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(32[13:44])
    inverter_U753 \inverter_chain_320..inv  (.\notGate[319]_keep (notGate_319), 
            .\notGate[320] (notGate_320)) /* synthesis syn_module_defined=1 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(32[13:44])
    inverter_U754 \inverter_chain_31..inv  (.\notGate[30]_keep (notGate_30), 
            .\notGate[31] (notGate_31)) /* synthesis syn_module_defined=1 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(32[13:44])
    inverter_U755 \inverter_chain_319..inv  (.\notGate[318]_keep (notGate_318), 
            .\notGate[319] (notGate_319)) /* synthesis syn_module_defined=1 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(32[13:44])
    inverter_U756 \inverter_chain_318..inv  (.\notGate[317]_keep (notGate_317), 
            .\notGate[318] (notGate_318)) /* synthesis syn_module_defined=1 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(32[13:44])
    inverter_U757 \inverter_chain_317..inv  (.\notGate[316]_keep (notGate_316), 
            .\notGate[317] (notGate_317)) /* synthesis syn_module_defined=1 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(32[13:44])
    inverter_U758 \inverter_chain_316..inv  (.\notGate[315]_keep (notGate_315), 
            .\notGate[316] (notGate_316)) /* synthesis syn_module_defined=1 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(32[13:44])
    inverter_U759 \inverter_chain_315..inv  (.\notGate[314]_keep (notGate_314), 
            .\notGate[315] (notGate_315)) /* synthesis syn_module_defined=1 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(32[13:44])
    inverter_U760 \inverter_chain_314..inv  (.\notGate[313]_keep (notGate_313), 
            .\notGate[314] (notGate_314)) /* synthesis syn_module_defined=1 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(32[13:44])
    inverter_U761 \inverter_chain_313..inv  (.\notGate[312]_keep (notGate_312), 
            .\notGate[313] (notGate_313)) /* synthesis syn_module_defined=1 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(32[13:44])
    inverter_U762 \inverter_chain_312..inv  (.\notGate[311]_keep (notGate_311), 
            .\notGate[312] (notGate_312)) /* synthesis syn_module_defined=1 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(32[13:44])
    inverter_U763 \inverter_chain_311..inv  (.\notGate[310]_keep (notGate_310), 
            .\notGate[311] (notGate_311)) /* synthesis syn_module_defined=1 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(32[13:44])
    inverter_U764 \inverter_chain_310..inv  (.\notGate[309]_keep (notGate_309), 
            .\notGate[310] (notGate_310)) /* synthesis syn_module_defined=1 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(32[13:44])
    inverter_U765 \inverter_chain_30..inv  (.\notGate[29]_keep (notGate_29), 
            .\notGate[30] (notGate_30)) /* synthesis syn_module_defined=1 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(32[13:44])
    inverter_U766 \inverter_chain_309..inv  (.\notGate[308]_keep (notGate_308), 
            .\notGate[309] (notGate_309)) /* synthesis syn_module_defined=1 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(32[13:44])
    inverter_U767 \inverter_chain_308..inv  (.\notGate[307]_keep (notGate_307), 
            .\notGate[308] (notGate_308)) /* synthesis syn_module_defined=1 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(32[13:44])
    inverter_U768 \inverter_chain_307..inv  (.\notGate[306]_keep (notGate_306), 
            .\notGate[307] (notGate_307)) /* synthesis syn_module_defined=1 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(32[13:44])
    inverter_U769 \inverter_chain_306..inv  (.\notGate[305]_keep (notGate_305), 
            .\notGate[306] (notGate_306)) /* synthesis syn_module_defined=1 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(32[13:44])
    inverter_U770 \inverter_chain_305..inv  (.\notGate[304]_keep (notGate_304), 
            .\notGate[305] (notGate_305)) /* synthesis syn_module_defined=1 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(32[13:44])
    inverter_U771 \inverter_chain_304..inv  (.\notGate[303]_keep (notGate_303), 
            .\notGate[304] (notGate_304)) /* synthesis syn_module_defined=1 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(32[13:44])
    inverter_U772 \inverter_chain_303..inv  (.\notGate[302]_keep (notGate_302), 
            .\notGate[303] (notGate_303)) /* synthesis syn_module_defined=1 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(32[13:44])
    inverter_U773 \inverter_chain_302..inv  (.\notGate[301]_keep (notGate_301), 
            .\notGate[302] (notGate_302)) /* synthesis syn_module_defined=1 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(32[13:44])
    inverter_U774 \inverter_chain_301..inv  (.\notGate[300]_keep (notGate_300), 
            .\notGate[301] (notGate_301)) /* synthesis syn_module_defined=1 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(32[13:44])
    inverter_U775 \inverter_chain_300..inv  (.\notGate[299]_keep (notGate_299), 
            .\notGate[300] (notGate_300)) /* synthesis syn_module_defined=1 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(32[13:44])
    inverter_U776 \inverter_chain_2..inv  (.\notGate[1]_keep (notGate_1), 
            .\notGate[2] (notGate_2)) /* synthesis syn_module_defined=1 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(32[13:44])
    inverter_U777 \inverter_chain_29..inv  (.\notGate[28]_keep (notGate_28), 
            .\notGate[29] (notGate_29)) /* synthesis syn_module_defined=1 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(32[13:44])
    inverter_U778 \inverter_chain_299..inv  (.\notGate[298]_keep (notGate_298), 
            .\notGate[299] (notGate_299)) /* synthesis syn_module_defined=1 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(32[13:44])
    inverter_U779 \inverter_chain_298..inv  (.\notGate[297]_keep (notGate_297), 
            .\notGate[298] (notGate_298)) /* synthesis syn_module_defined=1 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(32[13:44])
    inverter_U780 \inverter_chain_297..inv  (.\notGate[296]_keep (notGate_296), 
            .\notGate[297] (notGate_297)) /* synthesis syn_module_defined=1 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(32[13:44])
    inverter_U781 \inverter_chain_296..inv  (.\notGate[295]_keep (notGate_295), 
            .\notGate[296] (notGate_296)) /* synthesis syn_module_defined=1 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(32[13:44])
    inverter_U782 \inverter_chain_295..inv  (.\notGate[294]_keep (notGate_294), 
            .\notGate[295] (notGate_295)) /* synthesis syn_module_defined=1 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(32[13:44])
    inverter_U783 \inverter_chain_294..inv  (.\notGate[293]_keep (notGate_293), 
            .\notGate[294] (notGate_294)) /* synthesis syn_module_defined=1 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(32[13:44])
    inverter_U784 \inverter_chain_293..inv  (.\notGate[292]_keep (notGate_292), 
            .\notGate[293] (notGate_293)) /* synthesis syn_module_defined=1 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(32[13:44])
    inverter_U785 \inverter_chain_292..inv  (.\notGate[291]_keep (notGate_291), 
            .\notGate[292] (notGate_292)) /* synthesis syn_module_defined=1 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(32[13:44])
    inverter_U786 \inverter_chain_291..inv  (.\notGate[290]_keep (notGate_290), 
            .\notGate[291] (notGate_291)) /* synthesis syn_module_defined=1 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(32[13:44])
    inverter_U787 \inverter_chain_290..inv  (.\notGate[289]_keep (notGate_289), 
            .\notGate[290] (notGate_290)) /* synthesis syn_module_defined=1 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(32[13:44])
    inverter_U788 \inverter_chain_28..inv  (.\notGate[27]_keep (notGate_27), 
            .\notGate[28] (notGate_28)) /* synthesis syn_module_defined=1 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(32[13:44])
    inverter_U789 \inverter_chain_289..inv  (.\notGate[288]_keep (notGate_288), 
            .\notGate[289] (notGate_289)) /* synthesis syn_module_defined=1 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(32[13:44])
    inverter_U790 \inverter_chain_288..inv  (.\notGate[287]_keep (notGate_287), 
            .\notGate[288] (notGate_288)) /* synthesis syn_module_defined=1 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(32[13:44])
    inverter_U791 \inverter_chain_287..inv  (.\notGate[286]_keep (notGate_286), 
            .\notGate[287] (notGate_287)) /* synthesis syn_module_defined=1 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(32[13:44])
    inverter_U792 \inverter_chain_286..inv  (.\notGate[285]_keep (notGate_285), 
            .\notGate[286] (notGate_286)) /* synthesis syn_module_defined=1 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(32[13:44])
    inverter_U793 \inverter_chain_285..inv  (.\notGate[284]_keep (notGate_284), 
            .\notGate[285] (notGate_285)) /* synthesis syn_module_defined=1 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(32[13:44])
    inverter_U794 \inverter_chain_284..inv  (.\notGate[283]_keep (notGate_283), 
            .\notGate[284] (notGate_284)) /* synthesis syn_module_defined=1 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(32[13:44])
    inverter_U795 \inverter_chain_283..inv  (.\notGate[282]_keep (notGate_282), 
            .\notGate[283] (notGate_283)) /* synthesis syn_module_defined=1 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(32[13:44])
    inverter_U796 \inverter_chain_282..inv  (.\notGate[281]_keep (notGate_281), 
            .\notGate[282] (notGate_282)) /* synthesis syn_module_defined=1 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(32[13:44])
    inverter_U797 \inverter_chain_281..inv  (.\notGate[280]_keep (notGate_280), 
            .\notGate[281] (notGate_281)) /* synthesis syn_module_defined=1 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(32[13:44])
    inverter_U798 \inverter_chain_280..inv  (.\notGate[279]_keep (notGate_279), 
            .\notGate[280] (notGate_280)) /* synthesis syn_module_defined=1 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(32[13:44])
    inverter_U799 \inverter_chain_27..inv  (.\notGate[26]_keep (notGate_26), 
            .\notGate[27] (notGate_27)) /* synthesis syn_module_defined=1 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(32[13:44])
    inverter_U800 \inverter_chain_279..inv  (.\notGate[278]_keep (notGate_278), 
            .\notGate[279] (notGate_279)) /* synthesis syn_module_defined=1 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(32[13:44])
    inverter_U801 \inverter_chain_278..inv  (.\notGate[277]_keep (notGate_277), 
            .\notGate[278] (notGate_278)) /* synthesis syn_module_defined=1 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(32[13:44])
    inverter_U802 \inverter_chain_277..inv  (.\notGate[276]_keep (notGate_276), 
            .\notGate[277] (notGate_277)) /* synthesis syn_module_defined=1 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(32[13:44])
    inverter_U803 \inverter_chain_276..inv  (.\notGate[275]_keep (notGate_275), 
            .\notGate[276] (notGate_276)) /* synthesis syn_module_defined=1 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(32[13:44])
    inverter_U804 \inverter_chain_275..inv  (.\notGate[274]_keep (notGate_274), 
            .\notGate[275] (notGate_275)) /* synthesis syn_module_defined=1 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(32[13:44])
    inverter_U805 \inverter_chain_274..inv  (.\notGate[273]_keep (notGate_273), 
            .\notGate[274] (notGate_274)) /* synthesis syn_module_defined=1 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(32[13:44])
    inverter_U806 \inverter_chain_273..inv  (.\notGate[272]_keep (notGate_272), 
            .\notGate[273] (notGate_273)) /* synthesis syn_module_defined=1 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(32[13:44])
    inverter_U807 \inverter_chain_272..inv  (.\notGate[271]_keep (notGate_271), 
            .\notGate[272] (notGate_272)) /* synthesis syn_module_defined=1 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(32[13:44])
    inverter_U808 \inverter_chain_271..inv  (.\notGate[270]_keep (notGate_270), 
            .\notGate[271] (notGate_271)) /* synthesis syn_module_defined=1 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(32[13:44])
    inverter_U809 \inverter_chain_270..inv  (.\notGate[269]_keep (notGate_269), 
            .\notGate[270] (notGate_270)) /* synthesis syn_module_defined=1 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(32[13:44])
    inverter_U810 \inverter_chain_26..inv  (.\notGate[25]_keep (notGate_25), 
            .\notGate[26] (notGate_26)) /* synthesis syn_module_defined=1 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(32[13:44])
    inverter_U811 \inverter_chain_269..inv  (.\notGate[268]_keep (notGate_268), 
            .\notGate[269] (notGate_269)) /* synthesis syn_module_defined=1 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(32[13:44])
    inverter_U812 \inverter_chain_268..inv  (.\notGate[267]_keep (notGate_267), 
            .\notGate[268] (notGate_268)) /* synthesis syn_module_defined=1 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(32[13:44])
    inverter_U813 \inverter_chain_267..inv  (.\notGate[266]_keep (notGate_266), 
            .\notGate[267] (notGate_267)) /* synthesis syn_module_defined=1 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(32[13:44])
    inverter_U814 \inverter_chain_266..inv  (.\notGate[265]_keep (notGate_265), 
            .\notGate[266] (notGate_266)) /* synthesis syn_module_defined=1 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(32[13:44])
    inverter_U815 \inverter_chain_265..inv  (.\notGate[264]_keep (notGate_264), 
            .\notGate[265] (notGate_265)) /* synthesis syn_module_defined=1 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(32[13:44])
    inverter_U816 \inverter_chain_264..inv  (.\notGate[263]_keep (notGate_263), 
            .\notGate[264] (notGate_264)) /* synthesis syn_module_defined=1 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(32[13:44])
    inverter_U817 \inverter_chain_263..inv  (.\notGate[262]_keep (notGate_262), 
            .\notGate[263] (notGate_263)) /* synthesis syn_module_defined=1 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(32[13:44])
    inverter_U818 \inverter_chain_262..inv  (.\notGate[261]_keep (notGate_261), 
            .\notGate[262] (notGate_262)) /* synthesis syn_module_defined=1 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(32[13:44])
    inverter_U819 \inverter_chain_261..inv  (.\notGate[260]_keep (notGate_260), 
            .\notGate[261] (notGate_261)) /* synthesis syn_module_defined=1 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(32[13:44])
    inverter_U820 \inverter_chain_260..inv  (.\notGate[259]_keep (notGate_259), 
            .\notGate[260] (notGate_260)) /* synthesis syn_module_defined=1 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(32[13:44])
    inverter_U821 \inverter_chain_25..inv  (.\notGate[24]_keep (notGate_24), 
            .\notGate[25] (notGate_25)) /* synthesis syn_module_defined=1 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(32[13:44])
    inverter_U822 \inverter_chain_259..inv  (.\notGate[258]_keep (notGate_258), 
            .\notGate[259] (notGate_259)) /* synthesis syn_module_defined=1 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(32[13:44])
    inverter_U823 \inverter_chain_258..inv  (.\notGate[257]_keep (notGate_257), 
            .\notGate[258] (notGate_258)) /* synthesis syn_module_defined=1 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(32[13:44])
    inverter_U824 \inverter_chain_257..inv  (.\notGate[256]_keep (notGate_256), 
            .\notGate[257] (notGate_257)) /* synthesis syn_module_defined=1 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(32[13:44])
    inverter_U825 \inverter_chain_256..inv  (.\notGate[255]_keep (notGate_255), 
            .\notGate[256] (notGate_256)) /* synthesis syn_module_defined=1 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(32[13:44])
    inverter_U826 \inverter_chain_255..inv  (.\notGate[254]_keep (notGate_254), 
            .\notGate[255] (notGate_255)) /* synthesis syn_module_defined=1 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(32[13:44])
    inverter_U827 \inverter_chain_254..inv  (.\notGate[253]_keep (notGate_253), 
            .\notGate[254] (notGate_254)) /* synthesis syn_module_defined=1 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(32[13:44])
    inverter_U828 \inverter_chain_253..inv  (.\notGate[252]_keep (notGate_252), 
            .\notGate[253] (notGate_253)) /* synthesis syn_module_defined=1 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(32[13:44])
    inverter_U829 \inverter_chain_252..inv  (.\notGate[251]_keep (notGate_251), 
            .\notGate[252] (notGate_252)) /* synthesis syn_module_defined=1 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(32[13:44])
    inverter_U830 \inverter_chain_251..inv  (.\notGate[250]_keep (notGate_250), 
            .\notGate[251] (notGate_251)) /* synthesis syn_module_defined=1 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(32[13:44])
    inverter_U831 \inverter_chain_250..inv  (.\notGate[249]_keep (notGate_249), 
            .\notGate[250] (notGate_250)) /* synthesis syn_module_defined=1 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(32[13:44])
    inverter_U832 \inverter_chain_24..inv  (.\notGate[23]_keep (notGate_23), 
            .\notGate[24] (notGate_24)) /* synthesis syn_module_defined=1 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(32[13:44])
    inverter_U833 \inverter_chain_249..inv  (.\notGate[248]_keep (notGate_248), 
            .\notGate[249] (notGate_249)) /* synthesis syn_module_defined=1 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(32[13:44])
    inverter_U834 \inverter_chain_248..inv  (.\notGate[247]_keep (notGate_247), 
            .\notGate[248] (notGate_248)) /* synthesis syn_module_defined=1 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(32[13:44])
    inverter_U835 \inverter_chain_247..inv  (.\notGate[246]_keep (notGate_246), 
            .\notGate[247] (notGate_247)) /* synthesis syn_module_defined=1 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(32[13:44])
    inverter_U836 \inverter_chain_246..inv  (.\notGate[245]_keep (notGate_245), 
            .\notGate[246] (notGate_246)) /* synthesis syn_module_defined=1 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(32[13:44])
    inverter_U837 \inverter_chain_245..inv  (.\notGate[244]_keep (notGate_244), 
            .\notGate[245] (notGate_245)) /* synthesis syn_module_defined=1 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(32[13:44])
    inverter_U838 \inverter_chain_244..inv  (.\notGate[243]_keep (notGate_243), 
            .\notGate[244] (notGate_244)) /* synthesis syn_module_defined=1 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(32[13:44])
    inverter_U839 \inverter_chain_243..inv  (.\notGate[242]_keep (notGate_242), 
            .\notGate[243] (notGate_243)) /* synthesis syn_module_defined=1 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(32[13:44])
    inverter_U840 \inverter_chain_242..inv  (.\notGate[241]_keep (notGate_241), 
            .\notGate[242] (notGate_242)) /* synthesis syn_module_defined=1 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(32[13:44])
    inverter_U841 \inverter_chain_241..inv  (.\notGate[240]_keep (notGate_240), 
            .\notGate[241] (notGate_241)) /* synthesis syn_module_defined=1 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(32[13:44])
    inverter_U842 \inverter_chain_240..inv  (.\notGate[239]_keep (notGate_239), 
            .\notGate[240] (notGate_240)) /* synthesis syn_module_defined=1 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(32[13:44])
    inverter_U843 \inverter_chain_23..inv  (.\notGate[22]_keep (notGate_22), 
            .\notGate[23] (notGate_23)) /* synthesis syn_module_defined=1 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(32[13:44])
    inverter_U844 \inverter_chain_239..inv  (.\notGate[238]_keep (notGate_238), 
            .\notGate[239] (notGate_239)) /* synthesis syn_module_defined=1 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(32[13:44])
    inverter_U845 \inverter_chain_238..inv  (.\notGate[237]_keep (notGate_237), 
            .\notGate[238] (notGate_238)) /* synthesis syn_module_defined=1 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(32[13:44])
    inverter_U846 \inverter_chain_237..inv  (.\notGate[236]_keep (notGate_236), 
            .\notGate[237] (notGate_237)) /* synthesis syn_module_defined=1 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(32[13:44])
    inverter_U847 \inverter_chain_236..inv  (.\notGate[235]_keep (notGate_235), 
            .\notGate[236] (notGate_236)) /* synthesis syn_module_defined=1 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(32[13:44])
    inverter_U848 \inverter_chain_235..inv  (.\notGate[234]_keep (notGate_234), 
            .\notGate[235] (notGate_235)) /* synthesis syn_module_defined=1 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(32[13:44])
    inverter_U849 \inverter_chain_234..inv  (.\notGate[233]_keep (notGate_233), 
            .\notGate[234] (notGate_234)) /* synthesis syn_module_defined=1 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(32[13:44])
    inverter_U850 \inverter_chain_233..inv  (.\notGate[232]_keep (notGate_232), 
            .\notGate[233] (notGate_233)) /* synthesis syn_module_defined=1 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(32[13:44])
    inverter_U851 \inverter_chain_232..inv  (.\notGate[231]_keep (notGate_231), 
            .\notGate[232] (notGate_232)) /* synthesis syn_module_defined=1 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(32[13:44])
    inverter_U852 \inverter_chain_231..inv  (.\notGate[230]_keep (notGate_230), 
            .\notGate[231] (notGate_231)) /* synthesis syn_module_defined=1 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(32[13:44])
    inverter_U853 \inverter_chain_230..inv  (.\notGate[229]_keep (notGate_229), 
            .\notGate[230] (notGate_230)) /* synthesis syn_module_defined=1 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(32[13:44])
    inverter_U854 \inverter_chain_22..inv  (.\notGate[21]_keep (notGate_21), 
            .\notGate[22] (notGate_22)) /* synthesis syn_module_defined=1 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(32[13:44])
    inverter_U855 \inverter_chain_229..inv  (.\notGate[228]_keep (notGate_228), 
            .\notGate[229] (notGate_229)) /* synthesis syn_module_defined=1 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(32[13:44])
    inverter_U856 \inverter_chain_228..inv  (.\notGate[227]_keep (notGate_227), 
            .\notGate[228] (notGate_228)) /* synthesis syn_module_defined=1 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(32[13:44])
    inverter_U857 \inverter_chain_227..inv  (.\notGate[226]_keep (notGate_226), 
            .\notGate[227] (notGate_227)) /* synthesis syn_module_defined=1 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(32[13:44])
    inverter_U858 \inverter_chain_226..inv  (.\notGate[225]_keep (notGate_225), 
            .\notGate[226] (notGate_226)) /* synthesis syn_module_defined=1 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(32[13:44])
    inverter_U859 \inverter_chain_225..inv  (.\notGate[224]_keep (notGate_224), 
            .\notGate[225] (notGate_225)) /* synthesis syn_module_defined=1 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(32[13:44])
    inverter_U860 \inverter_chain_224..inv  (.\notGate[223]_keep (notGate_223), 
            .\notGate[224] (notGate_224)) /* synthesis syn_module_defined=1 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(32[13:44])
    inverter_U861 \inverter_chain_223..inv  (.\notGate[222]_keep (notGate_222), 
            .\notGate[223] (notGate_223)) /* synthesis syn_module_defined=1 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(32[13:44])
    inverter_U862 \inverter_chain_222..inv  (.\notGate[221]_keep (notGate_221), 
            .\notGate[222] (notGate_222)) /* synthesis syn_module_defined=1 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(32[13:44])
    inverter_U863 \inverter_chain_221..inv  (.\notGate[220]_keep (notGate_220), 
            .\notGate[221] (notGate_221)) /* synthesis syn_module_defined=1 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(32[13:44])
    inverter_U864 \inverter_chain_220..inv  (.\notGate[219]_keep (notGate_219), 
            .\notGate[220] (notGate_220)) /* synthesis syn_module_defined=1 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(32[13:44])
    inverter_U865 \inverter_chain_21..inv  (.\notGate[20]_keep (notGate_20), 
            .\notGate[21] (notGate_21)) /* synthesis syn_module_defined=1 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(32[13:44])
    inverter_U866 \inverter_chain_219..inv  (.\notGate[218]_keep (notGate_218), 
            .\notGate[219] (notGate_219)) /* synthesis syn_module_defined=1 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(32[13:44])
    inverter_U867 \inverter_chain_218..inv  (.\notGate[217]_keep (notGate_217), 
            .\notGate[218] (notGate_218)) /* synthesis syn_module_defined=1 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(32[13:44])
    inverter_U868 \inverter_chain_217..inv  (.\notGate[216]_keep (notGate_216), 
            .\notGate[217] (notGate_217)) /* synthesis syn_module_defined=1 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(32[13:44])
    inverter_U869 \inverter_chain_216..inv  (.\notGate[215]_keep (notGate_215), 
            .\notGate[216] (notGate_216)) /* synthesis syn_module_defined=1 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(32[13:44])
    inverter_U870 \inverter_chain_215..inv  (.\notGate[214]_keep (notGate_214), 
            .\notGate[215] (notGate_215)) /* synthesis syn_module_defined=1 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(32[13:44])
    inverter_U871 \inverter_chain_214..inv  (.\notGate[213]_keep (notGate_213), 
            .\notGate[214] (notGate_214)) /* synthesis syn_module_defined=1 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(32[13:44])
    inverter_U872 \inverter_chain_213..inv  (.\notGate[212]_keep (notGate_212), 
            .\notGate[213] (notGate_213)) /* synthesis syn_module_defined=1 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(32[13:44])
    inverter_U873 \inverter_chain_212..inv  (.\notGate[211]_keep (notGate_211), 
            .\notGate[212] (notGate_212)) /* synthesis syn_module_defined=1 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(32[13:44])
    inverter_U874 \inverter_chain_211..inv  (.\notGate[210]_keep (notGate_210), 
            .\notGate[211] (notGate_211)) /* synthesis syn_module_defined=1 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(32[13:44])
    inverter_U875 \inverter_chain_210..inv  (.\notGate[209]_keep (notGate_209), 
            .\notGate[210] (notGate_210)) /* synthesis syn_module_defined=1 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(32[13:44])
    inverter_U876 \inverter_chain_20..inv  (.\notGate[19]_keep (notGate_19), 
            .\notGate[20] (notGate_20)) /* synthesis syn_module_defined=1 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(32[13:44])
    inverter_U877 \inverter_chain_209..inv  (.\notGate[208]_keep (notGate_208), 
            .\notGate[209] (notGate_209)) /* synthesis syn_module_defined=1 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(32[13:44])
    inverter_U878 \inverter_chain_208..inv  (.\notGate[207]_keep (notGate_207), 
            .\notGate[208] (notGate_208)) /* synthesis syn_module_defined=1 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(32[13:44])
    inverter_U879 \inverter_chain_207..inv  (.\notGate[206]_keep (notGate_206), 
            .\notGate[207] (notGate_207)) /* synthesis syn_module_defined=1 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(32[13:44])
    inverter_U880 \inverter_chain_206..inv  (.\notGate[205]_keep (notGate_205), 
            .\notGate[206] (notGate_206)) /* synthesis syn_module_defined=1 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(32[13:44])
    inverter_U881 \inverter_chain_205..inv  (.\notGate[204]_keep (notGate_204), 
            .\notGate[205] (notGate_205)) /* synthesis syn_module_defined=1 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(32[13:44])
    inverter_U882 \inverter_chain_204..inv  (.\notGate[203]_keep (notGate_203), 
            .\notGate[204] (notGate_204)) /* synthesis syn_module_defined=1 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(32[13:44])
    inverter_U883 \inverter_chain_203..inv  (.\notGate[202]_keep (notGate_202), 
            .\notGate[203] (notGate_203)) /* synthesis syn_module_defined=1 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(32[13:44])
    inverter_U884 \inverter_chain_202..inv  (.\notGate[201]_keep (notGate_201), 
            .\notGate[202] (notGate_202)) /* synthesis syn_module_defined=1 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(32[13:44])
    inverter_U885 \inverter_chain_201..inv  (.\notGate[200]_keep (notGate_200), 
            .\notGate[201] (notGate_201)) /* synthesis syn_module_defined=1 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(32[13:44])
    inverter_U886 \inverter_chain_200..inv  (.\notGate[199]_keep (notGate_199), 
            .\notGate[200] (notGate_200)) /* synthesis syn_module_defined=1 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(32[13:44])
    inverter_U887 \inverter_chain_1..inv  (.\notGate[0]_keep (notGate_0), 
            .\notGate[1] (notGate_1)) /* synthesis syn_module_defined=1 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(32[13:44])
    inverter_U888 \inverter_chain_19..inv  (.\notGate[18]_keep (notGate_18), 
            .\notGate[19] (notGate_19)) /* synthesis syn_module_defined=1 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(32[13:44])
    inverter_U889 \inverter_chain_199..inv  (.\notGate[198]_keep (notGate_198), 
            .\notGate[199] (notGate_199)) /* synthesis syn_module_defined=1 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(32[13:44])
    inverter_U890 \inverter_chain_198..inv  (.\notGate[197]_keep (notGate_197), 
            .\notGate[198] (notGate_198)) /* synthesis syn_module_defined=1 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(32[13:44])
    inverter_U891 \inverter_chain_197..inv  (.\notGate[196]_keep (notGate_196), 
            .\notGate[197] (notGate_197)) /* synthesis syn_module_defined=1 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(32[13:44])
    inverter_U892 \inverter_chain_196..inv  (.\notGate[195]_keep (notGate_195), 
            .\notGate[196] (notGate_196)) /* synthesis syn_module_defined=1 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(32[13:44])
    inverter_U893 \inverter_chain_195..inv  (.\notGate[194]_keep (notGate_194), 
            .\notGate[195] (notGate_195)) /* synthesis syn_module_defined=1 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(32[13:44])
    inverter_U894 \inverter_chain_194..inv  (.\notGate[193]_keep (notGate_193), 
            .\notGate[194] (notGate_194)) /* synthesis syn_module_defined=1 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(32[13:44])
    inverter_U895 \inverter_chain_193..inv  (.\notGate[192]_keep (notGate_192), 
            .\notGate[193] (notGate_193)) /* synthesis syn_module_defined=1 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(32[13:44])
    inverter_U896 \inverter_chain_192..inv  (.\notGate[191]_keep (notGate_191), 
            .\notGate[192] (notGate_192)) /* synthesis syn_module_defined=1 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(32[13:44])
    inverter_U897 \inverter_chain_191..inv  (.\notGate[190]_keep (notGate_190), 
            .\notGate[191] (notGate_191)) /* synthesis syn_module_defined=1 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(32[13:44])
    inverter_U898 \inverter_chain_190..inv  (.\notGate[189]_keep (notGate_189), 
            .\notGate[190] (notGate_190)) /* synthesis syn_module_defined=1 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(32[13:44])
    inverter_U899 \inverter_chain_18..inv  (.\notGate[17]_keep (notGate_17), 
            .\notGate[18] (notGate_18)) /* synthesis syn_module_defined=1 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(32[13:44])
    inverter_U900 \inverter_chain_189..inv  (.\notGate[188]_keep (notGate_188), 
            .\notGate[189] (notGate_189)) /* synthesis syn_module_defined=1 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(32[13:44])
    inverter_U901 \inverter_chain_188..inv  (.\notGate[187]_keep (notGate_187), 
            .\notGate[188] (notGate_188)) /* synthesis syn_module_defined=1 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(32[13:44])
    inverter_U902 \inverter_chain_187..inv  (.\notGate[186]_keep (notGate_186), 
            .\notGate[187] (notGate_187)) /* synthesis syn_module_defined=1 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(32[13:44])
    inverter_U903 \inverter_chain_186..inv  (.\notGate[185]_keep (notGate_185), 
            .\notGate[186] (notGate_186)) /* synthesis syn_module_defined=1 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(32[13:44])
    inverter_U904 \inverter_chain_185..inv  (.\notGate[184]_keep (notGate_184), 
            .\notGate[185] (notGate_185)) /* synthesis syn_module_defined=1 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(32[13:44])
    inverter_U905 \inverter_chain_184..inv  (.\notGate[183]_keep (notGate_183), 
            .\notGate[184] (notGate_184)) /* synthesis syn_module_defined=1 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(32[13:44])
    inverter_U906 \inverter_chain_183..inv  (.\notGate[182]_keep (notGate_182), 
            .\notGate[183] (notGate_183)) /* synthesis syn_module_defined=1 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(32[13:44])
    inverter_U907 \inverter_chain_182..inv  (.\notGate[181]_keep (notGate_181), 
            .\notGate[182] (notGate_182)) /* synthesis syn_module_defined=1 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(32[13:44])
    inverter_U908 \inverter_chain_181..inv  (.\notGate[180]_keep (notGate_180), 
            .\notGate[181] (notGate_181)) /* synthesis syn_module_defined=1 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(32[13:44])
    inverter_U909 \inverter_chain_180..inv  (.\notGate[179]_keep (notGate_179), 
            .\notGate[180] (notGate_180)) /* synthesis syn_module_defined=1 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(32[13:44])
    inverter_U910 \inverter_chain_17..inv  (.\notGate[16]_keep (notGate_16), 
            .\notGate[17] (notGate_17)) /* synthesis syn_module_defined=1 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(32[13:44])
    inverter_U911 \inverter_chain_179..inv  (.\notGate[178]_keep (notGate_178), 
            .\notGate[179] (notGate_179)) /* synthesis syn_module_defined=1 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(32[13:44])
    inverter_U912 \inverter_chain_178..inv  (.\notGate[177]_keep (notGate_177), 
            .\notGate[178] (notGate_178)) /* synthesis syn_module_defined=1 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(32[13:44])
    inverter_U913 \inverter_chain_177..inv  (.\notGate[176]_keep (notGate_176), 
            .\notGate[177] (notGate_177)) /* synthesis syn_module_defined=1 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(32[13:44])
    inverter_U914 \inverter_chain_176..inv  (.\notGate[175]_keep (notGate_175), 
            .\notGate[176] (notGate_176)) /* synthesis syn_module_defined=1 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(32[13:44])
    inverter_U915 \inverter_chain_175..inv  (.\notGate[174]_keep (notGate_174), 
            .\notGate[175] (notGate_175)) /* synthesis syn_module_defined=1 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(32[13:44])
    inverter_U916 \inverter_chain_174..inv  (.\notGate[173]_keep (notGate_173), 
            .\notGate[174] (notGate_174)) /* synthesis syn_module_defined=1 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(32[13:44])
    inverter_U917 \inverter_chain_173..inv  (.\notGate[172]_keep (notGate_172), 
            .\notGate[173] (notGate_173)) /* synthesis syn_module_defined=1 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(32[13:44])
    inverter_U918 \inverter_chain_172..inv  (.\notGate[171]_keep (notGate_171), 
            .\notGate[172] (notGate_172)) /* synthesis syn_module_defined=1 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(32[13:44])
    inverter_U919 \inverter_chain_171..inv  (.\notGate[170]_keep (notGate_170), 
            .\notGate[171] (notGate_171)) /* synthesis syn_module_defined=1 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(32[13:44])
    inverter_U920 \inverter_chain_170..inv  (.\notGate[169]_keep (notGate_169), 
            .\notGate[170] (notGate_170)) /* synthesis syn_module_defined=1 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(32[13:44])
    inverter_U921 \inverter_chain_16..inv  (.\notGate[15]_keep (notGate_15), 
            .\notGate[16] (notGate_16)) /* synthesis syn_module_defined=1 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(32[13:44])
    inverter_U922 \inverter_chain_169..inv  (.\notGate[168]_keep (notGate_168), 
            .\notGate[169] (notGate_169)) /* synthesis syn_module_defined=1 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(32[13:44])
    inverter_U923 \inverter_chain_168..inv  (.\notGate[167]_keep (notGate_167), 
            .\notGate[168] (notGate_168)) /* synthesis syn_module_defined=1 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(32[13:44])
    inverter_U924 \inverter_chain_167..inv  (.\notGate[166]_keep (notGate_166), 
            .\notGate[167] (notGate_167)) /* synthesis syn_module_defined=1 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(32[13:44])
    inverter_U925 \inverter_chain_166..inv  (.\notGate[165]_keep (notGate_165), 
            .\notGate[166] (notGate_166)) /* synthesis syn_module_defined=1 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(32[13:44])
    inverter_U926 \inverter_chain_165..inv  (.\notGate[164]_keep (notGate_164), 
            .\notGate[165] (notGate_165)) /* synthesis syn_module_defined=1 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(32[13:44])
    inverter_U927 \inverter_chain_164..inv  (.\notGate[163]_keep (notGate_163), 
            .\notGate[164] (notGate_164)) /* synthesis syn_module_defined=1 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(32[13:44])
    inverter_U928 \inverter_chain_163..inv  (.\notGate[162]_keep (notGate_162), 
            .\notGate[163] (notGate_163)) /* synthesis syn_module_defined=1 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(32[13:44])
    inverter_U929 \inverter_chain_162..inv  (.\notGate[161]_keep (notGate_161), 
            .\notGate[162] (notGate_162)) /* synthesis syn_module_defined=1 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(32[13:44])
    inverter_U930 \inverter_chain_161..inv  (.\notGate[160]_keep (notGate_160), 
            .\notGate[161] (notGate_161)) /* synthesis syn_module_defined=1 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(32[13:44])
    inverter_U931 \inverter_chain_160..inv  (.\notGate[159]_keep (notGate_159), 
            .\notGate[160] (notGate_160)) /* synthesis syn_module_defined=1 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(32[13:44])
    inverter_U932 \inverter_chain_15..inv  (.\notGate[14]_keep (notGate_14), 
            .\notGate[15] (notGate_15)) /* synthesis syn_module_defined=1 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(32[13:44])
    inverter_U933 \inverter_chain_159..inv  (.\notGate[158]_keep (notGate_158), 
            .\notGate[159] (notGate_159)) /* synthesis syn_module_defined=1 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(32[13:44])
    inverter_U934 \inverter_chain_158..inv  (.\notGate[157]_keep (notGate_157), 
            .\notGate[158] (notGate_158)) /* synthesis syn_module_defined=1 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(32[13:44])
    inverter_U935 \inverter_chain_157..inv  (.\notGate[156]_keep (notGate_156), 
            .\notGate[157] (notGate_157)) /* synthesis syn_module_defined=1 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(32[13:44])
    inverter_U936 \inverter_chain_156..inv  (.\notGate[155]_keep (notGate_155), 
            .\notGate[156] (notGate_156)) /* synthesis syn_module_defined=1 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(32[13:44])
    inverter_U937 \inverter_chain_155..inv  (.\notGate[154]_keep (notGate_154), 
            .\notGate[155] (notGate_155)) /* synthesis syn_module_defined=1 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(32[13:44])
    inverter_U938 \inverter_chain_154..inv  (.\notGate[153]_keep (notGate_153), 
            .\notGate[154] (notGate_154)) /* synthesis syn_module_defined=1 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(32[13:44])
    inverter_U939 \inverter_chain_153..inv  (.\notGate[152]_keep (notGate_152), 
            .\notGate[153] (notGate_153)) /* synthesis syn_module_defined=1 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(32[13:44])
    inverter_U940 \inverter_chain_152..inv  (.\notGate[151]_keep (notGate_151), 
            .\notGate[152] (notGate_152)) /* synthesis syn_module_defined=1 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(32[13:44])
    inverter_U941 \inverter_chain_151..inv  (.\notGate[150]_keep (notGate_150), 
            .\notGate[151] (notGate_151)) /* synthesis syn_module_defined=1 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(32[13:44])
    inverter_U942 \inverter_chain_150..inv  (.\notGate[149]_keep (notGate_149), 
            .\notGate[150] (notGate_150)) /* synthesis syn_module_defined=1 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(32[13:44])
    inverter_U943 \inverter_chain_14..inv  (.\notGate[13]_keep (notGate_13), 
            .\notGate[14] (notGate_14)) /* synthesis syn_module_defined=1 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(32[13:44])
    inverter_U944 \inverter_chain_149..inv  (.\notGate[148]_keep (notGate_148), 
            .\notGate[149] (notGate_149)) /* synthesis syn_module_defined=1 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(32[13:44])
    inverter_U945 \inverter_chain_148..inv  (.\notGate[147]_keep (notGate_147), 
            .\notGate[148] (notGate_148)) /* synthesis syn_module_defined=1 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(32[13:44])
    inverter_U946 \inverter_chain_147..inv  (.\notGate[146]_keep (notGate_146), 
            .\notGate[147] (notGate_147)) /* synthesis syn_module_defined=1 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(32[13:44])
    inverter_U947 \inverter_chain_146..inv  (.\notGate[145]_keep (notGate_145), 
            .\notGate[146] (notGate_146)) /* synthesis syn_module_defined=1 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(32[13:44])
    inverter_U948 \inverter_chain_145..inv  (.\notGate[144]_keep (notGate_144), 
            .\notGate[145] (notGate_145)) /* synthesis syn_module_defined=1 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(32[13:44])
    inverter_U949 \inverter_chain_144..inv  (.\notGate[143]_keep (notGate_143), 
            .\notGate[144] (notGate_144)) /* synthesis syn_module_defined=1 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(32[13:44])
    inverter_U950 \inverter_chain_143..inv  (.\notGate[142]_keep (notGate_142), 
            .\notGate[143] (notGate_143)) /* synthesis syn_module_defined=1 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(32[13:44])
    inverter_U951 \inverter_chain_142..inv  (.\notGate[141]_keep (notGate_141), 
            .\notGate[142] (notGate_142)) /* synthesis syn_module_defined=1 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(32[13:44])
    inverter_U952 \inverter_chain_141..inv  (.\notGate[140]_keep (notGate_140), 
            .\notGate[141] (notGate_141)) /* synthesis syn_module_defined=1 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(32[13:44])
    inverter_U953 \inverter_chain_140..inv  (.\notGate[139]_keep (notGate_139), 
            .\notGate[140] (notGate_140)) /* synthesis syn_module_defined=1 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(32[13:44])
    inverter_U954 \inverter_chain_13..inv  (.\notGate[12]_keep (notGate_12), 
            .\notGate[13] (notGate_13)) /* synthesis syn_module_defined=1 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(32[13:44])
    inverter_U955 \inverter_chain_139..inv  (.\notGate[138]_keep (notGate_138), 
            .\notGate[139] (notGate_139)) /* synthesis syn_module_defined=1 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(32[13:44])
    inverter_U956 \inverter_chain_138..inv  (.\notGate[137]_keep (notGate_137), 
            .\notGate[138] (notGate_138)) /* synthesis syn_module_defined=1 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(32[13:44])
    inverter_U957 \inverter_chain_137..inv  (.\notGate[136]_keep (notGate_136), 
            .\notGate[137] (notGate_137)) /* synthesis syn_module_defined=1 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(32[13:44])
    inverter_U958 \inverter_chain_136..inv  (.\notGate[135]_keep (notGate_135), 
            .\notGate[136] (notGate_136)) /* synthesis syn_module_defined=1 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(32[13:44])
    inverter_U959 \inverter_chain_135..inv  (.\notGate[134]_keep (notGate_134), 
            .\notGate[135] (notGate_135)) /* synthesis syn_module_defined=1 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(32[13:44])
    inverter_U960 \inverter_chain_134..inv  (.\notGate[133]_keep (notGate_133), 
            .\notGate[134] (notGate_134)) /* synthesis syn_module_defined=1 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(32[13:44])
    inverter_U961 \inverter_chain_133..inv  (.\notGate[132]_keep (notGate_132), 
            .\notGate[133] (notGate_133)) /* synthesis syn_module_defined=1 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(32[13:44])
    inverter_U962 \inverter_chain_132..inv  (.\notGate[131]_keep (notGate_131), 
            .\notGate[132] (notGate_132)) /* synthesis syn_module_defined=1 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(32[13:44])
    inverter_U963 \inverter_chain_131..inv  (.\notGate[130]_keep (notGate_130), 
            .\notGate[131] (notGate_131)) /* synthesis syn_module_defined=1 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(32[13:44])
    inverter_U964 \inverter_chain_130..inv  (.\notGate[129]_keep (notGate_129), 
            .\notGate[130] (notGate_130)) /* synthesis syn_module_defined=1 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(32[13:44])
    inverter_U965 \inverter_chain_12..inv  (.\notGate[11]_keep (notGate_11), 
            .\notGate[12] (notGate_12)) /* synthesis syn_module_defined=1 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(32[13:44])
    inverter_U966 \inverter_chain_129..inv  (.\notGate[128]_keep (notGate_128), 
            .\notGate[129] (notGate_129)) /* synthesis syn_module_defined=1 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(32[13:44])
    inverter_U967 \inverter_chain_128..inv  (.\notGate[127]_keep (notGate_127), 
            .\notGate[128] (notGate_128)) /* synthesis syn_module_defined=1 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(32[13:44])
    inverter_U968 \inverter_chain_127..inv  (.\notGate[126]_keep (notGate_126), 
            .\notGate[127] (notGate_127)) /* synthesis syn_module_defined=1 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(32[13:44])
    inverter_U969 \inverter_chain_126..inv  (.\notGate[125]_keep (notGate_125), 
            .\notGate[126] (notGate_126)) /* synthesis syn_module_defined=1 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(32[13:44])
    inverter_U970 \inverter_chain_125..inv  (.\notGate[124]_keep (notGate_124), 
            .\notGate[125] (notGate_125)) /* synthesis syn_module_defined=1 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(32[13:44])
    inverter_U971 \inverter_chain_124..inv  (.\notGate[123]_keep (notGate_123), 
            .\notGate[124] (notGate_124)) /* synthesis syn_module_defined=1 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(32[13:44])
    inverter_U972 \inverter_chain_123..inv  (.\notGate[122]_keep (notGate_122), 
            .\notGate[123] (notGate_123)) /* synthesis syn_module_defined=1 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(32[13:44])
    inverter_U973 \inverter_chain_122..inv  (.\notGate[121]_keep (notGate_121), 
            .\notGate[122] (notGate_122)) /* synthesis syn_module_defined=1 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(32[13:44])
    inverter_U974 \inverter_chain_121..inv  (.\notGate[120]_keep (notGate_120), 
            .\notGate[121] (notGate_121)) /* synthesis syn_module_defined=1 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(32[13:44])
    inverter_U975 \inverter_chain_120..inv  (.\notGate[119]_keep (notGate_119), 
            .\notGate[120] (notGate_120)) /* synthesis syn_module_defined=1 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(32[13:44])
    inverter_U976 \inverter_chain_11..inv  (.\notGate[10]_keep (notGate_10), 
            .\notGate[11] (notGate_11)) /* synthesis syn_module_defined=1 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(32[13:44])
    inverter_U977 \inverter_chain_119..inv  (.\notGate[118]_keep (notGate_118), 
            .\notGate[119] (notGate_119)) /* synthesis syn_module_defined=1 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(32[13:44])
    inverter_U978 \inverter_chain_118..inv  (.\notGate[117]_keep (notGate_117), 
            .\notGate[118] (notGate_118)) /* synthesis syn_module_defined=1 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(32[13:44])
    inverter_U979 \inverter_chain_117..inv  (.\notGate[116]_keep (notGate_116), 
            .\notGate[117] (notGate_117)) /* synthesis syn_module_defined=1 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(32[13:44])
    inverter_U980 \inverter_chain_116..inv  (.\notGate[115]_keep (notGate_115), 
            .\notGate[116] (notGate_116)) /* synthesis syn_module_defined=1 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(32[13:44])
    inverter_U981 \inverter_chain_115..inv  (.\notGate[114]_keep (notGate_114), 
            .\notGate[115] (notGate_115)) /* synthesis syn_module_defined=1 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(32[13:44])
    inverter_U982 \inverter_chain_114..inv  (.\notGate[113]_keep (notGate_113), 
            .\notGate[114] (notGate_114)) /* synthesis syn_module_defined=1 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(32[13:44])
    inverter_U983 \inverter_chain_113..inv  (.\notGate[112]_keep (notGate_112), 
            .\notGate[113] (notGate_113)) /* synthesis syn_module_defined=1 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(32[13:44])
    inverter_U984 \inverter_chain_112..inv  (.\notGate[111]_keep (notGate_111), 
            .\notGate[112] (notGate_112)) /* synthesis syn_module_defined=1 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(32[13:44])
    inverter_U985 \inverter_chain_111..inv  (.\notGate[110]_keep (notGate_110), 
            .\notGate[111] (notGate_111)) /* synthesis syn_module_defined=1 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(32[13:44])
    inverter_U986 \inverter_chain_110..inv  (.\notGate[109]_keep (notGate_109), 
            .\notGate[110] (notGate_110)) /* synthesis syn_module_defined=1 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(32[13:44])
    inverter_U987 \inverter_chain_10..inv  (.\notGate[9]_keep (notGate_9), 
            .\notGate[10] (notGate_10)) /* synthesis syn_module_defined=1 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(32[13:44])
    inverter_U988 \inverter_chain_109..inv  (.\notGate[108]_keep (notGate_108), 
            .\notGate[109] (notGate_109)) /* synthesis syn_module_defined=1 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(32[13:44])
    inverter_U989 \inverter_chain_108..inv  (.\notGate[107]_keep (notGate_107), 
            .\notGate[108] (notGate_108)) /* synthesis syn_module_defined=1 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(32[13:44])
    inverter_U990 \inverter_chain_107..inv  (.\notGate[106]_keep (notGate_106), 
            .\notGate[107] (notGate_107)) /* synthesis syn_module_defined=1 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(32[13:44])
    inverter_U991 \inverter_chain_106..inv  (.\notGate[105]_keep (notGate_105), 
            .\notGate[106] (notGate_106)) /* synthesis syn_module_defined=1 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(32[13:44])
    inverter_U992 \inverter_chain_105..inv  (.\notGate[104]_keep (notGate_104), 
            .\notGate[105] (notGate_105)) /* synthesis syn_module_defined=1 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(32[13:44])
    inverter_U993 \inverter_chain_104..inv  (.\notGate[103]_keep (notGate_103), 
            .\notGate[104] (notGate_104)) /* synthesis syn_module_defined=1 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(32[13:44])
    inverter_U994 \inverter_chain_103..inv  (.\notGate[102]_keep (notGate_102), 
            .\notGate[103] (notGate_103)) /* synthesis syn_module_defined=1 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(32[13:44])
    inverter_U995 \inverter_chain_102..inv  (.\notGate[101]_keep (notGate_101), 
            .\notGate[102] (notGate_102)) /* synthesis syn_module_defined=1 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(32[13:44])
    inverter_U996 \inverter_chain_101..inv  (.\notGate[100]_keep (notGate_100), 
            .\notGate[101] (notGate_101)) /* synthesis syn_module_defined=1 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(32[13:44])
    inverter_U997 \inverter_chain_100..inv  (.\notGate[99]_keep (notGate_99), 
            .\notGate[100] (notGate_100)) /* synthesis syn_module_defined=1 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(32[13:44])
    inverter_U998 \inverter_chain_1000..inv  (.\notGate[999]_keep (notGate_999), 
            .\notGate[1000] (notGate_1000)) /* synthesis syn_module_defined=1 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(32[13:44])
    
endmodule
//
// Verilog Description of module inverter
//

module inverter (\notGate[8]_keep , \notGate[9] ) /* synthesis syn_module_defined=1 */ ;
    input \notGate[8]_keep ;
    output \notGate[9] ;
    
    wire \notGate[8]_keep  /* synthesis alspreserve=1 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(25[15:22])
    
    LUT4 I1 (.A(\notGate[8]_keep ), .B(\notGate[8]_keep ), .C(\notGate[8]_keep ), 
         .D(\notGate[8]_keep ), .Z(\notGate[9] )) /* synthesis syn_instantiated=1, lut_function=((!D !C !B !A)+(!D !C !B A)+(!D !C B !A)+(!D !C B A)+(!D C !B !A)+(!D C !B A)+(!D C B !A)+(!D C B A)), LSE_LINE_FILE_ID=3, LSE_LCOL=13, LSE_RCOL=44, LSE_LLINE=32, LSE_RLINE=32 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(11[2:53])
    defparam I1.init = 16'b0000000011111111;
    
endmodule
//
// Verilog Description of module inverter_U0
//

module inverter_U0 (\notGate[98]_keep , \notGate[99] ) /* synthesis syn_module_defined=1 */ ;
    input \notGate[98]_keep ;
    output \notGate[99] ;
    
    wire \notGate[98]_keep  /* synthesis alspreserve=1 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(25[15:22])
    
    LUT4 I1 (.A(\notGate[98]_keep ), .B(\notGate[98]_keep ), .C(\notGate[98]_keep ), 
         .D(\notGate[98]_keep ), .Z(\notGate[99] )) /* synthesis syn_instantiated=1, lut_function=((!D !C !B !A)+(!D !C !B A)+(!D !C B !A)+(!D !C B A)+(!D C !B !A)+(!D C !B A)+(!D C B !A)+(!D C B A)), LSE_LINE_FILE_ID=3, LSE_LCOL=13, LSE_RCOL=44, LSE_LLINE=32, LSE_RLINE=32 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(11[2:53])
    defparam I1.init = 16'b0000000011111111;
    
endmodule
//
// Verilog Description of module inverter_U1
//

module inverter_U1 (\notGate[998]_keep , \notGate[999] ) /* synthesis syn_module_defined=1 */ ;
    input \notGate[998]_keep ;
    output \notGate[999] ;
    
    wire \notGate[998]_keep  /* synthesis alspreserve=1 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(25[15:22])
    
    LUT4 I1 (.A(\notGate[998]_keep ), .B(\notGate[998]_keep ), .C(\notGate[998]_keep ), 
         .D(\notGate[998]_keep ), .Z(\notGate[999] )) /* synthesis syn_instantiated=1, lut_function=((!D !C !B !A)+(!D !C !B A)+(!D !C B !A)+(!D !C B A)+(!D C !B !A)+(!D C !B A)+(!D C B !A)+(!D C B A)), LSE_LINE_FILE_ID=3, LSE_LCOL=13, LSE_RCOL=44, LSE_LLINE=32, LSE_RLINE=32 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(11[2:53])
    defparam I1.init = 16'b0000000011111111;
    
endmodule
//
// Verilog Description of module inverter_U2
//

module inverter_U2 (\notGate[997]_keep , \notGate[998] ) /* synthesis syn_module_defined=1 */ ;
    input \notGate[997]_keep ;
    output \notGate[998] ;
    
    wire \notGate[997]_keep  /* synthesis alspreserve=1 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(25[15:22])
    
    LUT4 I1 (.A(\notGate[997]_keep ), .B(\notGate[997]_keep ), .C(\notGate[997]_keep ), 
         .D(\notGate[997]_keep ), .Z(\notGate[998] )) /* synthesis syn_instantiated=1, lut_function=((!D !C !B !A)+(!D !C !B A)+(!D !C B !A)+(!D !C B A)+(!D C !B !A)+(!D C !B A)+(!D C B !A)+(!D C B A)), LSE_LINE_FILE_ID=3, LSE_LCOL=13, LSE_RCOL=44, LSE_LLINE=32, LSE_RLINE=32 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(11[2:53])
    defparam I1.init = 16'b0000000011111111;
    
endmodule
//
// Verilog Description of module inverter_U3
//

module inverter_U3 (\notGate[996]_keep , \notGate[997] ) /* synthesis syn_module_defined=1 */ ;
    input \notGate[996]_keep ;
    output \notGate[997] ;
    
    wire \notGate[996]_keep  /* synthesis alspreserve=1 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(25[15:22])
    
    LUT4 I1 (.A(\notGate[996]_keep ), .B(\notGate[996]_keep ), .C(\notGate[996]_keep ), 
         .D(\notGate[996]_keep ), .Z(\notGate[997] )) /* synthesis syn_instantiated=1, lut_function=((!D !C !B !A)+(!D !C !B A)+(!D !C B !A)+(!D !C B A)+(!D C !B !A)+(!D C !B A)+(!D C B !A)+(!D C B A)), LSE_LINE_FILE_ID=3, LSE_LCOL=13, LSE_RCOL=44, LSE_LLINE=32, LSE_RLINE=32 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(11[2:53])
    defparam I1.init = 16'b0000000011111111;
    
endmodule
//
// Verilog Description of module inverter_U4
//

module inverter_U4 (\notGate[995]_keep , \notGate[996] ) /* synthesis syn_module_defined=1 */ ;
    input \notGate[995]_keep ;
    output \notGate[996] ;
    
    wire \notGate[995]_keep  /* synthesis alspreserve=1 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(25[15:22])
    
    LUT4 I1 (.A(\notGate[995]_keep ), .B(\notGate[995]_keep ), .C(\notGate[995]_keep ), 
         .D(\notGate[995]_keep ), .Z(\notGate[996] )) /* synthesis syn_instantiated=1, lut_function=((!D !C !B !A)+(!D !C !B A)+(!D !C B !A)+(!D !C B A)+(!D C !B !A)+(!D C !B A)+(!D C B !A)+(!D C B A)), LSE_LINE_FILE_ID=3, LSE_LCOL=13, LSE_RCOL=44, LSE_LLINE=32, LSE_RLINE=32 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(11[2:53])
    defparam I1.init = 16'b0000000011111111;
    
endmodule
//
// Verilog Description of module inverter_U5
//

module inverter_U5 (\notGate[994]_keep , \notGate[995] ) /* synthesis syn_module_defined=1 */ ;
    input \notGate[994]_keep ;
    output \notGate[995] ;
    
    wire \notGate[994]_keep  /* synthesis alspreserve=1 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(25[15:22])
    
    LUT4 I1 (.A(\notGate[994]_keep ), .B(\notGate[994]_keep ), .C(\notGate[994]_keep ), 
         .D(\notGate[994]_keep ), .Z(\notGate[995] )) /* synthesis syn_instantiated=1, lut_function=((!D !C !B !A)+(!D !C !B A)+(!D !C B !A)+(!D !C B A)+(!D C !B !A)+(!D C !B A)+(!D C B !A)+(!D C B A)), LSE_LINE_FILE_ID=3, LSE_LCOL=13, LSE_RCOL=44, LSE_LLINE=32, LSE_RLINE=32 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(11[2:53])
    defparam I1.init = 16'b0000000011111111;
    
endmodule
//
// Verilog Description of module inverter_U6
//

module inverter_U6 (\notGate[993]_keep , \notGate[994] ) /* synthesis syn_module_defined=1 */ ;
    input \notGate[993]_keep ;
    output \notGate[994] ;
    
    wire \notGate[993]_keep  /* synthesis alspreserve=1 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(25[15:22])
    
    LUT4 I1 (.A(\notGate[993]_keep ), .B(\notGate[993]_keep ), .C(\notGate[993]_keep ), 
         .D(\notGate[993]_keep ), .Z(\notGate[994] )) /* synthesis syn_instantiated=1, lut_function=((!D !C !B !A)+(!D !C !B A)+(!D !C B !A)+(!D !C B A)+(!D C !B !A)+(!D C !B A)+(!D C B !A)+(!D C B A)), LSE_LINE_FILE_ID=3, LSE_LCOL=13, LSE_RCOL=44, LSE_LLINE=32, LSE_RLINE=32 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(11[2:53])
    defparam I1.init = 16'b0000000011111111;
    
endmodule
//
// Verilog Description of module inverter_U7
//

module inverter_U7 (\notGate[992]_keep , \notGate[993] ) /* synthesis syn_module_defined=1 */ ;
    input \notGate[992]_keep ;
    output \notGate[993] ;
    
    wire \notGate[992]_keep  /* synthesis alspreserve=1 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(25[15:22])
    
    LUT4 I1 (.A(\notGate[992]_keep ), .B(\notGate[992]_keep ), .C(\notGate[992]_keep ), 
         .D(\notGate[992]_keep ), .Z(\notGate[993] )) /* synthesis syn_instantiated=1, lut_function=((!D !C !B !A)+(!D !C !B A)+(!D !C B !A)+(!D !C B A)+(!D C !B !A)+(!D C !B A)+(!D C B !A)+(!D C B A)), LSE_LINE_FILE_ID=3, LSE_LCOL=13, LSE_RCOL=44, LSE_LLINE=32, LSE_RLINE=32 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(11[2:53])
    defparam I1.init = 16'b0000000011111111;
    
endmodule
//
// Verilog Description of module inverter_U8
//

module inverter_U8 (\notGate[991]_keep , \notGate[992] ) /* synthesis syn_module_defined=1 */ ;
    input \notGate[991]_keep ;
    output \notGate[992] ;
    
    wire \notGate[991]_keep  /* synthesis alspreserve=1 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(25[15:22])
    
    LUT4 I1 (.A(\notGate[991]_keep ), .B(\notGate[991]_keep ), .C(\notGate[991]_keep ), 
         .D(\notGate[991]_keep ), .Z(\notGate[992] )) /* synthesis syn_instantiated=1, lut_function=((!D !C !B !A)+(!D !C !B A)+(!D !C B !A)+(!D !C B A)+(!D C !B !A)+(!D C !B A)+(!D C B !A)+(!D C B A)), LSE_LINE_FILE_ID=3, LSE_LCOL=13, LSE_RCOL=44, LSE_LLINE=32, LSE_RLINE=32 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(11[2:53])
    defparam I1.init = 16'b0000000011111111;
    
endmodule
//
// Verilog Description of module inverter_U9
//

module inverter_U9 (\notGate[990]_keep , \notGate[991] ) /* synthesis syn_module_defined=1 */ ;
    input \notGate[990]_keep ;
    output \notGate[991] ;
    
    wire \notGate[990]_keep  /* synthesis alspreserve=1 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(25[15:22])
    
    LUT4 I1 (.A(\notGate[990]_keep ), .B(\notGate[990]_keep ), .C(\notGate[990]_keep ), 
         .D(\notGate[990]_keep ), .Z(\notGate[991] )) /* synthesis syn_instantiated=1, lut_function=((!D !C !B !A)+(!D !C !B A)+(!D !C B !A)+(!D !C B A)+(!D C !B !A)+(!D C !B A)+(!D C B !A)+(!D C B A)), LSE_LINE_FILE_ID=3, LSE_LCOL=13, LSE_RCOL=44, LSE_LLINE=32, LSE_RLINE=32 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(11[2:53])
    defparam I1.init = 16'b0000000011111111;
    
endmodule
//
// Verilog Description of module inverter_U10
//

module inverter_U10 (\notGate[989]_keep , \notGate[990] ) /* synthesis syn_module_defined=1 */ ;
    input \notGate[989]_keep ;
    output \notGate[990] ;
    
    wire \notGate[989]_keep  /* synthesis alspreserve=1 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(25[15:22])
    
    LUT4 I1 (.A(\notGate[989]_keep ), .B(\notGate[989]_keep ), .C(\notGate[989]_keep ), 
         .D(\notGate[989]_keep ), .Z(\notGate[990] )) /* synthesis syn_instantiated=1, lut_function=((!D !C !B !A)+(!D !C !B A)+(!D !C B !A)+(!D !C B A)+(!D C !B !A)+(!D C !B A)+(!D C B !A)+(!D C B A)), LSE_LINE_FILE_ID=3, LSE_LCOL=13, LSE_RCOL=44, LSE_LLINE=32, LSE_RLINE=32 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(11[2:53])
    defparam I1.init = 16'b0000000011111111;
    
endmodule
//
// Verilog Description of module inverter_U11
//

module inverter_U11 (\notGate[97]_keep , \notGate[98] ) /* synthesis syn_module_defined=1 */ ;
    input \notGate[97]_keep ;
    output \notGate[98] ;
    
    wire \notGate[97]_keep  /* synthesis alspreserve=1 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(25[15:22])
    
    LUT4 I1 (.A(\notGate[97]_keep ), .B(\notGate[97]_keep ), .C(\notGate[97]_keep ), 
         .D(\notGate[97]_keep ), .Z(\notGate[98] )) /* synthesis syn_instantiated=1, lut_function=((!D !C !B !A)+(!D !C !B A)+(!D !C B !A)+(!D !C B A)+(!D C !B !A)+(!D C !B A)+(!D C B !A)+(!D C B A)), LSE_LINE_FILE_ID=3, LSE_LCOL=13, LSE_RCOL=44, LSE_LLINE=32, LSE_RLINE=32 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(11[2:53])
    defparam I1.init = 16'b0000000011111111;
    
endmodule
//
// Verilog Description of module inverter_U12
//

module inverter_U12 (\notGate[988]_keep , \notGate[989] ) /* synthesis syn_module_defined=1 */ ;
    input \notGate[988]_keep ;
    output \notGate[989] ;
    
    wire \notGate[988]_keep  /* synthesis alspreserve=1 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(25[15:22])
    
    LUT4 I1 (.A(\notGate[988]_keep ), .B(\notGate[988]_keep ), .C(\notGate[988]_keep ), 
         .D(\notGate[988]_keep ), .Z(\notGate[989] )) /* synthesis syn_instantiated=1, lut_function=((!D !C !B !A)+(!D !C !B A)+(!D !C B !A)+(!D !C B A)+(!D C !B !A)+(!D C !B A)+(!D C B !A)+(!D C B A)), LSE_LINE_FILE_ID=3, LSE_LCOL=13, LSE_RCOL=44, LSE_LLINE=32, LSE_RLINE=32 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(11[2:53])
    defparam I1.init = 16'b0000000011111111;
    
endmodule
//
// Verilog Description of module inverter_U13
//

module inverter_U13 (\notGate[987]_keep , \notGate[988] ) /* synthesis syn_module_defined=1 */ ;
    input \notGate[987]_keep ;
    output \notGate[988] ;
    
    wire \notGate[987]_keep  /* synthesis alspreserve=1 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(25[15:22])
    
    LUT4 I1 (.A(\notGate[987]_keep ), .B(\notGate[987]_keep ), .C(\notGate[987]_keep ), 
         .D(\notGate[987]_keep ), .Z(\notGate[988] )) /* synthesis syn_instantiated=1, lut_function=((!D !C !B !A)+(!D !C !B A)+(!D !C B !A)+(!D !C B A)+(!D C !B !A)+(!D C !B A)+(!D C B !A)+(!D C B A)), LSE_LINE_FILE_ID=3, LSE_LCOL=13, LSE_RCOL=44, LSE_LLINE=32, LSE_RLINE=32 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(11[2:53])
    defparam I1.init = 16'b0000000011111111;
    
endmodule
//
// Verilog Description of module inverter_U14
//

module inverter_U14 (\notGate[986]_keep , \notGate[987] ) /* synthesis syn_module_defined=1 */ ;
    input \notGate[986]_keep ;
    output \notGate[987] ;
    
    wire \notGate[986]_keep  /* synthesis alspreserve=1 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(25[15:22])
    
    LUT4 I1 (.A(\notGate[986]_keep ), .B(\notGate[986]_keep ), .C(\notGate[986]_keep ), 
         .D(\notGate[986]_keep ), .Z(\notGate[987] )) /* synthesis syn_instantiated=1, lut_function=((!D !C !B !A)+(!D !C !B A)+(!D !C B !A)+(!D !C B A)+(!D C !B !A)+(!D C !B A)+(!D C B !A)+(!D C B A)), LSE_LINE_FILE_ID=3, LSE_LCOL=13, LSE_RCOL=44, LSE_LLINE=32, LSE_RLINE=32 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(11[2:53])
    defparam I1.init = 16'b0000000011111111;
    
endmodule
//
// Verilog Description of module inverter_U15
//

module inverter_U15 (\notGate[985]_keep , \notGate[986] ) /* synthesis syn_module_defined=1 */ ;
    input \notGate[985]_keep ;
    output \notGate[986] ;
    
    wire \notGate[985]_keep  /* synthesis alspreserve=1 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(25[15:22])
    
    LUT4 I1 (.A(\notGate[985]_keep ), .B(\notGate[985]_keep ), .C(\notGate[985]_keep ), 
         .D(\notGate[985]_keep ), .Z(\notGate[986] )) /* synthesis syn_instantiated=1, lut_function=((!D !C !B !A)+(!D !C !B A)+(!D !C B !A)+(!D !C B A)+(!D C !B !A)+(!D C !B A)+(!D C B !A)+(!D C B A)), LSE_LINE_FILE_ID=3, LSE_LCOL=13, LSE_RCOL=44, LSE_LLINE=32, LSE_RLINE=32 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(11[2:53])
    defparam I1.init = 16'b0000000011111111;
    
endmodule
//
// Verilog Description of module inverter_U16
//

module inverter_U16 (\notGate[984]_keep , \notGate[985] ) /* synthesis syn_module_defined=1 */ ;
    input \notGate[984]_keep ;
    output \notGate[985] ;
    
    wire \notGate[984]_keep  /* synthesis alspreserve=1 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(25[15:22])
    
    LUT4 I1 (.A(\notGate[984]_keep ), .B(\notGate[984]_keep ), .C(\notGate[984]_keep ), 
         .D(\notGate[984]_keep ), .Z(\notGate[985] )) /* synthesis syn_instantiated=1, lut_function=((!D !C !B !A)+(!D !C !B A)+(!D !C B !A)+(!D !C B A)+(!D C !B !A)+(!D C !B A)+(!D C B !A)+(!D C B A)), LSE_LINE_FILE_ID=3, LSE_LCOL=13, LSE_RCOL=44, LSE_LLINE=32, LSE_RLINE=32 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(11[2:53])
    defparam I1.init = 16'b0000000011111111;
    
endmodule
//
// Verilog Description of module inverter_U17
//

module inverter_U17 (\notGate[983]_keep , \notGate[984] ) /* synthesis syn_module_defined=1 */ ;
    input \notGate[983]_keep ;
    output \notGate[984] ;
    
    wire \notGate[983]_keep  /* synthesis alspreserve=1 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(25[15:22])
    
    LUT4 I1 (.A(\notGate[983]_keep ), .B(\notGate[983]_keep ), .C(\notGate[983]_keep ), 
         .D(\notGate[983]_keep ), .Z(\notGate[984] )) /* synthesis syn_instantiated=1, lut_function=((!D !C !B !A)+(!D !C !B A)+(!D !C B !A)+(!D !C B A)+(!D C !B !A)+(!D C !B A)+(!D C B !A)+(!D C B A)), LSE_LINE_FILE_ID=3, LSE_LCOL=13, LSE_RCOL=44, LSE_LLINE=32, LSE_RLINE=32 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(11[2:53])
    defparam I1.init = 16'b0000000011111111;
    
endmodule
//
// Verilog Description of module inverter_U18
//

module inverter_U18 (\notGate[982]_keep , \notGate[983] ) /* synthesis syn_module_defined=1 */ ;
    input \notGate[982]_keep ;
    output \notGate[983] ;
    
    wire \notGate[982]_keep  /* synthesis alspreserve=1 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(25[15:22])
    
    LUT4 I1 (.A(\notGate[982]_keep ), .B(\notGate[982]_keep ), .C(\notGate[982]_keep ), 
         .D(\notGate[982]_keep ), .Z(\notGate[983] )) /* synthesis syn_instantiated=1, lut_function=((!D !C !B !A)+(!D !C !B A)+(!D !C B !A)+(!D !C B A)+(!D C !B !A)+(!D C !B A)+(!D C B !A)+(!D C B A)), LSE_LINE_FILE_ID=3, LSE_LCOL=13, LSE_RCOL=44, LSE_LLINE=32, LSE_RLINE=32 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(11[2:53])
    defparam I1.init = 16'b0000000011111111;
    
endmodule
//
// Verilog Description of module inverter_U19
//

module inverter_U19 (\notGate[981]_keep , \notGate[982] ) /* synthesis syn_module_defined=1 */ ;
    input \notGate[981]_keep ;
    output \notGate[982] ;
    
    wire \notGate[981]_keep  /* synthesis alspreserve=1 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(25[15:22])
    
    LUT4 I1 (.A(\notGate[981]_keep ), .B(\notGate[981]_keep ), .C(\notGate[981]_keep ), 
         .D(\notGate[981]_keep ), .Z(\notGate[982] )) /* synthesis syn_instantiated=1, lut_function=((!D !C !B !A)+(!D !C !B A)+(!D !C B !A)+(!D !C B A)+(!D C !B !A)+(!D C !B A)+(!D C B !A)+(!D C B A)), LSE_LINE_FILE_ID=3, LSE_LCOL=13, LSE_RCOL=44, LSE_LLINE=32, LSE_RLINE=32 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(11[2:53])
    defparam I1.init = 16'b0000000011111111;
    
endmodule
//
// Verilog Description of module inverter_U20
//

module inverter_U20 (\notGate[980]_keep , \notGate[981] ) /* synthesis syn_module_defined=1 */ ;
    input \notGate[980]_keep ;
    output \notGate[981] ;
    
    wire \notGate[980]_keep  /* synthesis alspreserve=1 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(25[15:22])
    
    LUT4 I1 (.A(\notGate[980]_keep ), .B(\notGate[980]_keep ), .C(\notGate[980]_keep ), 
         .D(\notGate[980]_keep ), .Z(\notGate[981] )) /* synthesis syn_instantiated=1, lut_function=((!D !C !B !A)+(!D !C !B A)+(!D !C B !A)+(!D !C B A)+(!D C !B !A)+(!D C !B A)+(!D C B !A)+(!D C B A)), LSE_LINE_FILE_ID=3, LSE_LCOL=13, LSE_RCOL=44, LSE_LLINE=32, LSE_RLINE=32 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(11[2:53])
    defparam I1.init = 16'b0000000011111111;
    
endmodule
//
// Verilog Description of module inverter_U21
//

module inverter_U21 (\notGate[979]_keep , \notGate[980] ) /* synthesis syn_module_defined=1 */ ;
    input \notGate[979]_keep ;
    output \notGate[980] ;
    
    wire \notGate[979]_keep  /* synthesis alspreserve=1 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(25[15:22])
    
    LUT4 I1 (.A(\notGate[979]_keep ), .B(\notGate[979]_keep ), .C(\notGate[979]_keep ), 
         .D(\notGate[979]_keep ), .Z(\notGate[980] )) /* synthesis syn_instantiated=1, lut_function=((!D !C !B !A)+(!D !C !B A)+(!D !C B !A)+(!D !C B A)+(!D C !B !A)+(!D C !B A)+(!D C B !A)+(!D C B A)), LSE_LINE_FILE_ID=3, LSE_LCOL=13, LSE_RCOL=44, LSE_LLINE=32, LSE_RLINE=32 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(11[2:53])
    defparam I1.init = 16'b0000000011111111;
    
endmodule
//
// Verilog Description of module inverter_U22
//

module inverter_U22 (\notGate[96]_keep , \notGate[97] ) /* synthesis syn_module_defined=1 */ ;
    input \notGate[96]_keep ;
    output \notGate[97] ;
    
    wire \notGate[96]_keep  /* synthesis alspreserve=1 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(25[15:22])
    
    LUT4 I1 (.A(\notGate[96]_keep ), .B(\notGate[96]_keep ), .C(\notGate[96]_keep ), 
         .D(\notGate[96]_keep ), .Z(\notGate[97] )) /* synthesis syn_instantiated=1, lut_function=((!D !C !B !A)+(!D !C !B A)+(!D !C B !A)+(!D !C B A)+(!D C !B !A)+(!D C !B A)+(!D C B !A)+(!D C B A)), LSE_LINE_FILE_ID=3, LSE_LCOL=13, LSE_RCOL=44, LSE_LLINE=32, LSE_RLINE=32 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(11[2:53])
    defparam I1.init = 16'b0000000011111111;
    
endmodule
//
// Verilog Description of module inverter_U23
//

module inverter_U23 (\notGate[978]_keep , \notGate[979] ) /* synthesis syn_module_defined=1 */ ;
    input \notGate[978]_keep ;
    output \notGate[979] ;
    
    wire \notGate[978]_keep  /* synthesis alspreserve=1 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(25[15:22])
    
    LUT4 I1 (.A(\notGate[978]_keep ), .B(\notGate[978]_keep ), .C(\notGate[978]_keep ), 
         .D(\notGate[978]_keep ), .Z(\notGate[979] )) /* synthesis syn_instantiated=1, lut_function=((!D !C !B !A)+(!D !C !B A)+(!D !C B !A)+(!D !C B A)+(!D C !B !A)+(!D C !B A)+(!D C B !A)+(!D C B A)), LSE_LINE_FILE_ID=3, LSE_LCOL=13, LSE_RCOL=44, LSE_LLINE=32, LSE_RLINE=32 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(11[2:53])
    defparam I1.init = 16'b0000000011111111;
    
endmodule
//
// Verilog Description of module inverter_U24
//

module inverter_U24 (\notGate[977]_keep , \notGate[978] ) /* synthesis syn_module_defined=1 */ ;
    input \notGate[977]_keep ;
    output \notGate[978] ;
    
    wire \notGate[977]_keep  /* synthesis alspreserve=1 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(25[15:22])
    
    LUT4 I1 (.A(\notGate[977]_keep ), .B(\notGate[977]_keep ), .C(\notGate[977]_keep ), 
         .D(\notGate[977]_keep ), .Z(\notGate[978] )) /* synthesis syn_instantiated=1, lut_function=((!D !C !B !A)+(!D !C !B A)+(!D !C B !A)+(!D !C B A)+(!D C !B !A)+(!D C !B A)+(!D C B !A)+(!D C B A)), LSE_LINE_FILE_ID=3, LSE_LCOL=13, LSE_RCOL=44, LSE_LLINE=32, LSE_RLINE=32 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(11[2:53])
    defparam I1.init = 16'b0000000011111111;
    
endmodule
//
// Verilog Description of module inverter_U25
//

module inverter_U25 (\notGate[976]_keep , \notGate[977] ) /* synthesis syn_module_defined=1 */ ;
    input \notGate[976]_keep ;
    output \notGate[977] ;
    
    wire \notGate[976]_keep  /* synthesis alspreserve=1 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(25[15:22])
    
    LUT4 I1 (.A(\notGate[976]_keep ), .B(\notGate[976]_keep ), .C(\notGate[976]_keep ), 
         .D(\notGate[976]_keep ), .Z(\notGate[977] )) /* synthesis syn_instantiated=1, lut_function=((!D !C !B !A)+(!D !C !B A)+(!D !C B !A)+(!D !C B A)+(!D C !B !A)+(!D C !B A)+(!D C B !A)+(!D C B A)), LSE_LINE_FILE_ID=3, LSE_LCOL=13, LSE_RCOL=44, LSE_LLINE=32, LSE_RLINE=32 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(11[2:53])
    defparam I1.init = 16'b0000000011111111;
    
endmodule
//
// Verilog Description of module inverter_U26
//

module inverter_U26 (\notGate[975]_keep , \notGate[976] ) /* synthesis syn_module_defined=1 */ ;
    input \notGate[975]_keep ;
    output \notGate[976] ;
    
    wire \notGate[975]_keep  /* synthesis alspreserve=1 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(25[15:22])
    
    LUT4 I1 (.A(\notGate[975]_keep ), .B(\notGate[975]_keep ), .C(\notGate[975]_keep ), 
         .D(\notGate[975]_keep ), .Z(\notGate[976] )) /* synthesis syn_instantiated=1, lut_function=((!D !C !B !A)+(!D !C !B A)+(!D !C B !A)+(!D !C B A)+(!D C !B !A)+(!D C !B A)+(!D C B !A)+(!D C B A)), LSE_LINE_FILE_ID=3, LSE_LCOL=13, LSE_RCOL=44, LSE_LLINE=32, LSE_RLINE=32 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(11[2:53])
    defparam I1.init = 16'b0000000011111111;
    
endmodule
//
// Verilog Description of module inverter_U27
//

module inverter_U27 (\notGate[974]_keep , \notGate[975] ) /* synthesis syn_module_defined=1 */ ;
    input \notGate[974]_keep ;
    output \notGate[975] ;
    
    wire \notGate[974]_keep  /* synthesis alspreserve=1 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(25[15:22])
    
    LUT4 I1 (.A(\notGate[974]_keep ), .B(\notGate[974]_keep ), .C(\notGate[974]_keep ), 
         .D(\notGate[974]_keep ), .Z(\notGate[975] )) /* synthesis syn_instantiated=1, lut_function=((!D !C !B !A)+(!D !C !B A)+(!D !C B !A)+(!D !C B A)+(!D C !B !A)+(!D C !B A)+(!D C B !A)+(!D C B A)), LSE_LINE_FILE_ID=3, LSE_LCOL=13, LSE_RCOL=44, LSE_LLINE=32, LSE_RLINE=32 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(11[2:53])
    defparam I1.init = 16'b0000000011111111;
    
endmodule
//
// Verilog Description of module inverter_U28
//

module inverter_U28 (\notGate[973]_keep , \notGate[974] ) /* synthesis syn_module_defined=1 */ ;
    input \notGate[973]_keep ;
    output \notGate[974] ;
    
    wire \notGate[973]_keep  /* synthesis alspreserve=1 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(25[15:22])
    
    LUT4 I1 (.A(\notGate[973]_keep ), .B(\notGate[973]_keep ), .C(\notGate[973]_keep ), 
         .D(\notGate[973]_keep ), .Z(\notGate[974] )) /* synthesis syn_instantiated=1, lut_function=((!D !C !B !A)+(!D !C !B A)+(!D !C B !A)+(!D !C B A)+(!D C !B !A)+(!D C !B A)+(!D C B !A)+(!D C B A)), LSE_LINE_FILE_ID=3, LSE_LCOL=13, LSE_RCOL=44, LSE_LLINE=32, LSE_RLINE=32 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(11[2:53])
    defparam I1.init = 16'b0000000011111111;
    
endmodule
//
// Verilog Description of module inverter_U29
//

module inverter_U29 (\notGate[972]_keep , \notGate[973] ) /* synthesis syn_module_defined=1 */ ;
    input \notGate[972]_keep ;
    output \notGate[973] ;
    
    wire \notGate[972]_keep  /* synthesis alspreserve=1 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(25[15:22])
    
    LUT4 I1 (.A(\notGate[972]_keep ), .B(\notGate[972]_keep ), .C(\notGate[972]_keep ), 
         .D(\notGate[972]_keep ), .Z(\notGate[973] )) /* synthesis syn_instantiated=1, lut_function=((!D !C !B !A)+(!D !C !B A)+(!D !C B !A)+(!D !C B A)+(!D C !B !A)+(!D C !B A)+(!D C B !A)+(!D C B A)), LSE_LINE_FILE_ID=3, LSE_LCOL=13, LSE_RCOL=44, LSE_LLINE=32, LSE_RLINE=32 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(11[2:53])
    defparam I1.init = 16'b0000000011111111;
    
endmodule
//
// Verilog Description of module inverter_U30
//

module inverter_U30 (\notGate[971]_keep , \notGate[972] ) /* synthesis syn_module_defined=1 */ ;
    input \notGate[971]_keep ;
    output \notGate[972] ;
    
    wire \notGate[971]_keep  /* synthesis alspreserve=1 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(25[15:22])
    
    LUT4 I1 (.A(\notGate[971]_keep ), .B(\notGate[971]_keep ), .C(\notGate[971]_keep ), 
         .D(\notGate[971]_keep ), .Z(\notGate[972] )) /* synthesis syn_instantiated=1, lut_function=((!D !C !B !A)+(!D !C !B A)+(!D !C B !A)+(!D !C B A)+(!D C !B !A)+(!D C !B A)+(!D C B !A)+(!D C B A)), LSE_LINE_FILE_ID=3, LSE_LCOL=13, LSE_RCOL=44, LSE_LLINE=32, LSE_RLINE=32 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(11[2:53])
    defparam I1.init = 16'b0000000011111111;
    
endmodule
//
// Verilog Description of module inverter_U31
//

module inverter_U31 (\notGate[970]_keep , \notGate[971] ) /* synthesis syn_module_defined=1 */ ;
    input \notGate[970]_keep ;
    output \notGate[971] ;
    
    wire \notGate[970]_keep  /* synthesis alspreserve=1 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(25[15:22])
    
    LUT4 I1 (.A(\notGate[970]_keep ), .B(\notGate[970]_keep ), .C(\notGate[970]_keep ), 
         .D(\notGate[970]_keep ), .Z(\notGate[971] )) /* synthesis syn_instantiated=1, lut_function=((!D !C !B !A)+(!D !C !B A)+(!D !C B !A)+(!D !C B A)+(!D C !B !A)+(!D C !B A)+(!D C B !A)+(!D C B A)), LSE_LINE_FILE_ID=3, LSE_LCOL=13, LSE_RCOL=44, LSE_LLINE=32, LSE_RLINE=32 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(11[2:53])
    defparam I1.init = 16'b0000000011111111;
    
endmodule
//
// Verilog Description of module inverter_U32
//

module inverter_U32 (\notGate[969]_keep , \notGate[970] ) /* synthesis syn_module_defined=1 */ ;
    input \notGate[969]_keep ;
    output \notGate[970] ;
    
    wire \notGate[969]_keep  /* synthesis alspreserve=1 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(25[15:22])
    
    LUT4 I1 (.A(\notGate[969]_keep ), .B(\notGate[969]_keep ), .C(\notGate[969]_keep ), 
         .D(\notGate[969]_keep ), .Z(\notGate[970] )) /* synthesis syn_instantiated=1, lut_function=((!D !C !B !A)+(!D !C !B A)+(!D !C B !A)+(!D !C B A)+(!D C !B !A)+(!D C !B A)+(!D C B !A)+(!D C B A)), LSE_LINE_FILE_ID=3, LSE_LCOL=13, LSE_RCOL=44, LSE_LLINE=32, LSE_RLINE=32 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(11[2:53])
    defparam I1.init = 16'b0000000011111111;
    
endmodule
//
// Verilog Description of module inverter_U33
//

module inverter_U33 (\notGate[95]_keep , \notGate[96] ) /* synthesis syn_module_defined=1 */ ;
    input \notGate[95]_keep ;
    output \notGate[96] ;
    
    wire \notGate[95]_keep  /* synthesis alspreserve=1 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(25[15:22])
    
    LUT4 I1 (.A(\notGate[95]_keep ), .B(\notGate[95]_keep ), .C(\notGate[95]_keep ), 
         .D(\notGate[95]_keep ), .Z(\notGate[96] )) /* synthesis syn_instantiated=1, lut_function=((!D !C !B !A)+(!D !C !B A)+(!D !C B !A)+(!D !C B A)+(!D C !B !A)+(!D C !B A)+(!D C B !A)+(!D C B A)), LSE_LINE_FILE_ID=3, LSE_LCOL=13, LSE_RCOL=44, LSE_LLINE=32, LSE_RLINE=32 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(11[2:53])
    defparam I1.init = 16'b0000000011111111;
    
endmodule
//
// Verilog Description of module inverter_U34
//

module inverter_U34 (\notGate[968]_keep , \notGate[969] ) /* synthesis syn_module_defined=1 */ ;
    input \notGate[968]_keep ;
    output \notGate[969] ;
    
    wire \notGate[968]_keep  /* synthesis alspreserve=1 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(25[15:22])
    
    LUT4 I1 (.A(\notGate[968]_keep ), .B(\notGate[968]_keep ), .C(\notGate[968]_keep ), 
         .D(\notGate[968]_keep ), .Z(\notGate[969] )) /* synthesis syn_instantiated=1, lut_function=((!D !C !B !A)+(!D !C !B A)+(!D !C B !A)+(!D !C B A)+(!D C !B !A)+(!D C !B A)+(!D C B !A)+(!D C B A)), LSE_LINE_FILE_ID=3, LSE_LCOL=13, LSE_RCOL=44, LSE_LLINE=32, LSE_RLINE=32 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(11[2:53])
    defparam I1.init = 16'b0000000011111111;
    
endmodule
//
// Verilog Description of module inverter_U35
//

module inverter_U35 (\notGate[967]_keep , \notGate[968] ) /* synthesis syn_module_defined=1 */ ;
    input \notGate[967]_keep ;
    output \notGate[968] ;
    
    wire \notGate[967]_keep  /* synthesis alspreserve=1 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(25[15:22])
    
    LUT4 I1 (.A(\notGate[967]_keep ), .B(\notGate[967]_keep ), .C(\notGate[967]_keep ), 
         .D(\notGate[967]_keep ), .Z(\notGate[968] )) /* synthesis syn_instantiated=1, lut_function=((!D !C !B !A)+(!D !C !B A)+(!D !C B !A)+(!D !C B A)+(!D C !B !A)+(!D C !B A)+(!D C B !A)+(!D C B A)), LSE_LINE_FILE_ID=3, LSE_LCOL=13, LSE_RCOL=44, LSE_LLINE=32, LSE_RLINE=32 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(11[2:53])
    defparam I1.init = 16'b0000000011111111;
    
endmodule
//
// Verilog Description of module inverter_U36
//

module inverter_U36 (\notGate[966]_keep , \notGate[967] ) /* synthesis syn_module_defined=1 */ ;
    input \notGate[966]_keep ;
    output \notGate[967] ;
    
    wire \notGate[966]_keep  /* synthesis alspreserve=1 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(25[15:22])
    
    LUT4 I1 (.A(\notGate[966]_keep ), .B(\notGate[966]_keep ), .C(\notGate[966]_keep ), 
         .D(\notGate[966]_keep ), .Z(\notGate[967] )) /* synthesis syn_instantiated=1, lut_function=((!D !C !B !A)+(!D !C !B A)+(!D !C B !A)+(!D !C B A)+(!D C !B !A)+(!D C !B A)+(!D C B !A)+(!D C B A)), LSE_LINE_FILE_ID=3, LSE_LCOL=13, LSE_RCOL=44, LSE_LLINE=32, LSE_RLINE=32 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(11[2:53])
    defparam I1.init = 16'b0000000011111111;
    
endmodule
//
// Verilog Description of module inverter_U37
//

module inverter_U37 (\notGate[965]_keep , \notGate[966] ) /* synthesis syn_module_defined=1 */ ;
    input \notGate[965]_keep ;
    output \notGate[966] ;
    
    wire \notGate[965]_keep  /* synthesis alspreserve=1 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(25[15:22])
    
    LUT4 I1 (.A(\notGate[965]_keep ), .B(\notGate[965]_keep ), .C(\notGate[965]_keep ), 
         .D(\notGate[965]_keep ), .Z(\notGate[966] )) /* synthesis syn_instantiated=1, lut_function=((!D !C !B !A)+(!D !C !B A)+(!D !C B !A)+(!D !C B A)+(!D C !B !A)+(!D C !B A)+(!D C B !A)+(!D C B A)), LSE_LINE_FILE_ID=3, LSE_LCOL=13, LSE_RCOL=44, LSE_LLINE=32, LSE_RLINE=32 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(11[2:53])
    defparam I1.init = 16'b0000000011111111;
    
endmodule
//
// Verilog Description of module inverter_U38
//

module inverter_U38 (\notGate[964]_keep , \notGate[965] ) /* synthesis syn_module_defined=1 */ ;
    input \notGate[964]_keep ;
    output \notGate[965] ;
    
    wire \notGate[964]_keep  /* synthesis alspreserve=1 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(25[15:22])
    
    LUT4 I1 (.A(\notGate[964]_keep ), .B(\notGate[964]_keep ), .C(\notGate[964]_keep ), 
         .D(\notGate[964]_keep ), .Z(\notGate[965] )) /* synthesis syn_instantiated=1, lut_function=((!D !C !B !A)+(!D !C !B A)+(!D !C B !A)+(!D !C B A)+(!D C !B !A)+(!D C !B A)+(!D C B !A)+(!D C B A)), LSE_LINE_FILE_ID=3, LSE_LCOL=13, LSE_RCOL=44, LSE_LLINE=32, LSE_RLINE=32 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(11[2:53])
    defparam I1.init = 16'b0000000011111111;
    
endmodule
//
// Verilog Description of module inverter_U39
//

module inverter_U39 (\notGate[963]_keep , \notGate[964] ) /* synthesis syn_module_defined=1 */ ;
    input \notGate[963]_keep ;
    output \notGate[964] ;
    
    wire \notGate[963]_keep  /* synthesis alspreserve=1 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(25[15:22])
    
    LUT4 I1 (.A(\notGate[963]_keep ), .B(\notGate[963]_keep ), .C(\notGate[963]_keep ), 
         .D(\notGate[963]_keep ), .Z(\notGate[964] )) /* synthesis syn_instantiated=1, lut_function=((!D !C !B !A)+(!D !C !B A)+(!D !C B !A)+(!D !C B A)+(!D C !B !A)+(!D C !B A)+(!D C B !A)+(!D C B A)), LSE_LINE_FILE_ID=3, LSE_LCOL=13, LSE_RCOL=44, LSE_LLINE=32, LSE_RLINE=32 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(11[2:53])
    defparam I1.init = 16'b0000000011111111;
    
endmodule
//
// Verilog Description of module inverter_U40
//

module inverter_U40 (\notGate[962]_keep , \notGate[963] ) /* synthesis syn_module_defined=1 */ ;
    input \notGate[962]_keep ;
    output \notGate[963] ;
    
    wire \notGate[962]_keep  /* synthesis alspreserve=1 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(25[15:22])
    
    LUT4 I1 (.A(\notGate[962]_keep ), .B(\notGate[962]_keep ), .C(\notGate[962]_keep ), 
         .D(\notGate[962]_keep ), .Z(\notGate[963] )) /* synthesis syn_instantiated=1, lut_function=((!D !C !B !A)+(!D !C !B A)+(!D !C B !A)+(!D !C B A)+(!D C !B !A)+(!D C !B A)+(!D C B !A)+(!D C B A)), LSE_LINE_FILE_ID=3, LSE_LCOL=13, LSE_RCOL=44, LSE_LLINE=32, LSE_RLINE=32 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(11[2:53])
    defparam I1.init = 16'b0000000011111111;
    
endmodule
//
// Verilog Description of module inverter_U41
//

module inverter_U41 (\notGate[961]_keep , \notGate[962] ) /* synthesis syn_module_defined=1 */ ;
    input \notGate[961]_keep ;
    output \notGate[962] ;
    
    wire \notGate[961]_keep  /* synthesis alspreserve=1 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(25[15:22])
    
    LUT4 I1 (.A(\notGate[961]_keep ), .B(\notGate[961]_keep ), .C(\notGate[961]_keep ), 
         .D(\notGate[961]_keep ), .Z(\notGate[962] )) /* synthesis syn_instantiated=1, lut_function=((!D !C !B !A)+(!D !C !B A)+(!D !C B !A)+(!D !C B A)+(!D C !B !A)+(!D C !B A)+(!D C B !A)+(!D C B A)), LSE_LINE_FILE_ID=3, LSE_LCOL=13, LSE_RCOL=44, LSE_LLINE=32, LSE_RLINE=32 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(11[2:53])
    defparam I1.init = 16'b0000000011111111;
    
endmodule
//
// Verilog Description of module inverter_U42
//

module inverter_U42 (\notGate[960]_keep , \notGate[961] ) /* synthesis syn_module_defined=1 */ ;
    input \notGate[960]_keep ;
    output \notGate[961] ;
    
    wire \notGate[960]_keep  /* synthesis alspreserve=1 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(25[15:22])
    
    LUT4 I1 (.A(\notGate[960]_keep ), .B(\notGate[960]_keep ), .C(\notGate[960]_keep ), 
         .D(\notGate[960]_keep ), .Z(\notGate[961] )) /* synthesis syn_instantiated=1, lut_function=((!D !C !B !A)+(!D !C !B A)+(!D !C B !A)+(!D !C B A)+(!D C !B !A)+(!D C !B A)+(!D C B !A)+(!D C B A)), LSE_LINE_FILE_ID=3, LSE_LCOL=13, LSE_RCOL=44, LSE_LLINE=32, LSE_RLINE=32 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(11[2:53])
    defparam I1.init = 16'b0000000011111111;
    
endmodule
//
// Verilog Description of module inverter_U43
//

module inverter_U43 (\notGate[959]_keep , \notGate[960] ) /* synthesis syn_module_defined=1 */ ;
    input \notGate[959]_keep ;
    output \notGate[960] ;
    
    wire \notGate[959]_keep  /* synthesis alspreserve=1 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(25[15:22])
    
    LUT4 I1 (.A(\notGate[959]_keep ), .B(\notGate[959]_keep ), .C(\notGate[959]_keep ), 
         .D(\notGate[959]_keep ), .Z(\notGate[960] )) /* synthesis syn_instantiated=1, lut_function=((!D !C !B !A)+(!D !C !B A)+(!D !C B !A)+(!D !C B A)+(!D C !B !A)+(!D C !B A)+(!D C B !A)+(!D C B A)), LSE_LINE_FILE_ID=3, LSE_LCOL=13, LSE_RCOL=44, LSE_LLINE=32, LSE_RLINE=32 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(11[2:53])
    defparam I1.init = 16'b0000000011111111;
    
endmodule
//
// Verilog Description of module inverter_U44
//

module inverter_U44 (\notGate[94]_keep , \notGate[95] ) /* synthesis syn_module_defined=1 */ ;
    input \notGate[94]_keep ;
    output \notGate[95] ;
    
    wire \notGate[94]_keep  /* synthesis alspreserve=1 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(25[15:22])
    
    LUT4 I1 (.A(\notGate[94]_keep ), .B(\notGate[94]_keep ), .C(\notGate[94]_keep ), 
         .D(\notGate[94]_keep ), .Z(\notGate[95] )) /* synthesis syn_instantiated=1, lut_function=((!D !C !B !A)+(!D !C !B A)+(!D !C B !A)+(!D !C B A)+(!D C !B !A)+(!D C !B A)+(!D C B !A)+(!D C B A)), LSE_LINE_FILE_ID=3, LSE_LCOL=13, LSE_RCOL=44, LSE_LLINE=32, LSE_RLINE=32 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(11[2:53])
    defparam I1.init = 16'b0000000011111111;
    
endmodule
//
// Verilog Description of module inverter_U45
//

module inverter_U45 (\notGate[958]_keep , \notGate[959] ) /* synthesis syn_module_defined=1 */ ;
    input \notGate[958]_keep ;
    output \notGate[959] ;
    
    wire \notGate[958]_keep  /* synthesis alspreserve=1 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(25[15:22])
    
    LUT4 I1 (.A(\notGate[958]_keep ), .B(\notGate[958]_keep ), .C(\notGate[958]_keep ), 
         .D(\notGate[958]_keep ), .Z(\notGate[959] )) /* synthesis syn_instantiated=1, lut_function=((!D !C !B !A)+(!D !C !B A)+(!D !C B !A)+(!D !C B A)+(!D C !B !A)+(!D C !B A)+(!D C B !A)+(!D C B A)), LSE_LINE_FILE_ID=3, LSE_LCOL=13, LSE_RCOL=44, LSE_LLINE=32, LSE_RLINE=32 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(11[2:53])
    defparam I1.init = 16'b0000000011111111;
    
endmodule
//
// Verilog Description of module inverter_U46
//

module inverter_U46 (\notGate[957]_keep , \notGate[958] ) /* synthesis syn_module_defined=1 */ ;
    input \notGate[957]_keep ;
    output \notGate[958] ;
    
    wire \notGate[957]_keep  /* synthesis alspreserve=1 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(25[15:22])
    
    LUT4 I1 (.A(\notGate[957]_keep ), .B(\notGate[957]_keep ), .C(\notGate[957]_keep ), 
         .D(\notGate[957]_keep ), .Z(\notGate[958] )) /* synthesis syn_instantiated=1, lut_function=((!D !C !B !A)+(!D !C !B A)+(!D !C B !A)+(!D !C B A)+(!D C !B !A)+(!D C !B A)+(!D C B !A)+(!D C B A)), LSE_LINE_FILE_ID=3, LSE_LCOL=13, LSE_RCOL=44, LSE_LLINE=32, LSE_RLINE=32 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(11[2:53])
    defparam I1.init = 16'b0000000011111111;
    
endmodule
//
// Verilog Description of module inverter_U47
//

module inverter_U47 (\notGate[956]_keep , \notGate[957] ) /* synthesis syn_module_defined=1 */ ;
    input \notGate[956]_keep ;
    output \notGate[957] ;
    
    wire \notGate[956]_keep  /* synthesis alspreserve=1 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(25[15:22])
    
    LUT4 I1 (.A(\notGate[956]_keep ), .B(\notGate[956]_keep ), .C(\notGate[956]_keep ), 
         .D(\notGate[956]_keep ), .Z(\notGate[957] )) /* synthesis syn_instantiated=1, lut_function=((!D !C !B !A)+(!D !C !B A)+(!D !C B !A)+(!D !C B A)+(!D C !B !A)+(!D C !B A)+(!D C B !A)+(!D C B A)), LSE_LINE_FILE_ID=3, LSE_LCOL=13, LSE_RCOL=44, LSE_LLINE=32, LSE_RLINE=32 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(11[2:53])
    defparam I1.init = 16'b0000000011111111;
    
endmodule
//
// Verilog Description of module inverter_U48
//

module inverter_U48 (\notGate[955]_keep , \notGate[956] ) /* synthesis syn_module_defined=1 */ ;
    input \notGate[955]_keep ;
    output \notGate[956] ;
    
    wire \notGate[955]_keep  /* synthesis alspreserve=1 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(25[15:22])
    
    LUT4 I1 (.A(\notGate[955]_keep ), .B(\notGate[955]_keep ), .C(\notGate[955]_keep ), 
         .D(\notGate[955]_keep ), .Z(\notGate[956] )) /* synthesis syn_instantiated=1, lut_function=((!D !C !B !A)+(!D !C !B A)+(!D !C B !A)+(!D !C B A)+(!D C !B !A)+(!D C !B A)+(!D C B !A)+(!D C B A)), LSE_LINE_FILE_ID=3, LSE_LCOL=13, LSE_RCOL=44, LSE_LLINE=32, LSE_RLINE=32 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(11[2:53])
    defparam I1.init = 16'b0000000011111111;
    
endmodule
//
// Verilog Description of module inverter_U49
//

module inverter_U49 (\notGate[954]_keep , \notGate[955] ) /* synthesis syn_module_defined=1 */ ;
    input \notGate[954]_keep ;
    output \notGate[955] ;
    
    wire \notGate[954]_keep  /* synthesis alspreserve=1 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(25[15:22])
    
    LUT4 I1 (.A(\notGate[954]_keep ), .B(\notGate[954]_keep ), .C(\notGate[954]_keep ), 
         .D(\notGate[954]_keep ), .Z(\notGate[955] )) /* synthesis syn_instantiated=1, lut_function=((!D !C !B !A)+(!D !C !B A)+(!D !C B !A)+(!D !C B A)+(!D C !B !A)+(!D C !B A)+(!D C B !A)+(!D C B A)), LSE_LINE_FILE_ID=3, LSE_LCOL=13, LSE_RCOL=44, LSE_LLINE=32, LSE_RLINE=32 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(11[2:53])
    defparam I1.init = 16'b0000000011111111;
    
endmodule
//
// Verilog Description of module inverter_U50
//

module inverter_U50 (\notGate[953]_keep , \notGate[954] ) /* synthesis syn_module_defined=1 */ ;
    input \notGate[953]_keep ;
    output \notGate[954] ;
    
    wire \notGate[953]_keep  /* synthesis alspreserve=1 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(25[15:22])
    
    LUT4 I1 (.A(\notGate[953]_keep ), .B(\notGate[953]_keep ), .C(\notGate[953]_keep ), 
         .D(\notGate[953]_keep ), .Z(\notGate[954] )) /* synthesis syn_instantiated=1, lut_function=((!D !C !B !A)+(!D !C !B A)+(!D !C B !A)+(!D !C B A)+(!D C !B !A)+(!D C !B A)+(!D C B !A)+(!D C B A)), LSE_LINE_FILE_ID=3, LSE_LCOL=13, LSE_RCOL=44, LSE_LLINE=32, LSE_RLINE=32 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(11[2:53])
    defparam I1.init = 16'b0000000011111111;
    
endmodule
//
// Verilog Description of module inverter_U51
//

module inverter_U51 (\notGate[952]_keep , \notGate[953] ) /* synthesis syn_module_defined=1 */ ;
    input \notGate[952]_keep ;
    output \notGate[953] ;
    
    wire \notGate[952]_keep  /* synthesis alspreserve=1 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(25[15:22])
    
    LUT4 I1 (.A(\notGate[952]_keep ), .B(\notGate[952]_keep ), .C(\notGate[952]_keep ), 
         .D(\notGate[952]_keep ), .Z(\notGate[953] )) /* synthesis syn_instantiated=1, lut_function=((!D !C !B !A)+(!D !C !B A)+(!D !C B !A)+(!D !C B A)+(!D C !B !A)+(!D C !B A)+(!D C B !A)+(!D C B A)), LSE_LINE_FILE_ID=3, LSE_LCOL=13, LSE_RCOL=44, LSE_LLINE=32, LSE_RLINE=32 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(11[2:53])
    defparam I1.init = 16'b0000000011111111;
    
endmodule
//
// Verilog Description of module inverter_U52
//

module inverter_U52 (\notGate[951]_keep , \notGate[952] ) /* synthesis syn_module_defined=1 */ ;
    input \notGate[951]_keep ;
    output \notGate[952] ;
    
    wire \notGate[951]_keep  /* synthesis alspreserve=1 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(25[15:22])
    
    LUT4 I1 (.A(\notGate[951]_keep ), .B(\notGate[951]_keep ), .C(\notGate[951]_keep ), 
         .D(\notGate[951]_keep ), .Z(\notGate[952] )) /* synthesis syn_instantiated=1, lut_function=((!D !C !B !A)+(!D !C !B A)+(!D !C B !A)+(!D !C B A)+(!D C !B !A)+(!D C !B A)+(!D C B !A)+(!D C B A)), LSE_LINE_FILE_ID=3, LSE_LCOL=13, LSE_RCOL=44, LSE_LLINE=32, LSE_RLINE=32 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(11[2:53])
    defparam I1.init = 16'b0000000011111111;
    
endmodule
//
// Verilog Description of module inverter_U53
//

module inverter_U53 (\notGate[950]_keep , \notGate[951] ) /* synthesis syn_module_defined=1 */ ;
    input \notGate[950]_keep ;
    output \notGate[951] ;
    
    wire \notGate[950]_keep  /* synthesis alspreserve=1 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(25[15:22])
    
    LUT4 I1 (.A(\notGate[950]_keep ), .B(\notGate[950]_keep ), .C(\notGate[950]_keep ), 
         .D(\notGate[950]_keep ), .Z(\notGate[951] )) /* synthesis syn_instantiated=1, lut_function=((!D !C !B !A)+(!D !C !B A)+(!D !C B !A)+(!D !C B A)+(!D C !B !A)+(!D C !B A)+(!D C B !A)+(!D C B A)), LSE_LINE_FILE_ID=3, LSE_LCOL=13, LSE_RCOL=44, LSE_LLINE=32, LSE_RLINE=32 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(11[2:53])
    defparam I1.init = 16'b0000000011111111;
    
endmodule
//
// Verilog Description of module inverter_U54
//

module inverter_U54 (\notGate[949]_keep , \notGate[950] ) /* synthesis syn_module_defined=1 */ ;
    input \notGate[949]_keep ;
    output \notGate[950] ;
    
    wire \notGate[949]_keep  /* synthesis alspreserve=1 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(25[15:22])
    
    LUT4 I1 (.A(\notGate[949]_keep ), .B(\notGate[949]_keep ), .C(\notGate[949]_keep ), 
         .D(\notGate[949]_keep ), .Z(\notGate[950] )) /* synthesis syn_instantiated=1, lut_function=((!D !C !B !A)+(!D !C !B A)+(!D !C B !A)+(!D !C B A)+(!D C !B !A)+(!D C !B A)+(!D C B !A)+(!D C B A)), LSE_LINE_FILE_ID=3, LSE_LCOL=13, LSE_RCOL=44, LSE_LLINE=32, LSE_RLINE=32 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(11[2:53])
    defparam I1.init = 16'b0000000011111111;
    
endmodule
//
// Verilog Description of module inverter_U55
//

module inverter_U55 (\notGate[93]_keep , \notGate[94] ) /* synthesis syn_module_defined=1 */ ;
    input \notGate[93]_keep ;
    output \notGate[94] ;
    
    wire \notGate[93]_keep  /* synthesis alspreserve=1 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(25[15:22])
    
    LUT4 I1 (.A(\notGate[93]_keep ), .B(\notGate[93]_keep ), .C(\notGate[93]_keep ), 
         .D(\notGate[93]_keep ), .Z(\notGate[94] )) /* synthesis syn_instantiated=1, lut_function=((!D !C !B !A)+(!D !C !B A)+(!D !C B !A)+(!D !C B A)+(!D C !B !A)+(!D C !B A)+(!D C B !A)+(!D C B A)), LSE_LINE_FILE_ID=3, LSE_LCOL=13, LSE_RCOL=44, LSE_LLINE=32, LSE_RLINE=32 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(11[2:53])
    defparam I1.init = 16'b0000000011111111;
    
endmodule
//
// Verilog Description of module inverter_U56
//

module inverter_U56 (\notGate[948]_keep , \notGate[949] ) /* synthesis syn_module_defined=1 */ ;
    input \notGate[948]_keep ;
    output \notGate[949] ;
    
    wire \notGate[948]_keep  /* synthesis alspreserve=1 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(25[15:22])
    
    LUT4 I1 (.A(\notGate[948]_keep ), .B(\notGate[948]_keep ), .C(\notGate[948]_keep ), 
         .D(\notGate[948]_keep ), .Z(\notGate[949] )) /* synthesis syn_instantiated=1, lut_function=((!D !C !B !A)+(!D !C !B A)+(!D !C B !A)+(!D !C B A)+(!D C !B !A)+(!D C !B A)+(!D C B !A)+(!D C B A)), LSE_LINE_FILE_ID=3, LSE_LCOL=13, LSE_RCOL=44, LSE_LLINE=32, LSE_RLINE=32 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(11[2:53])
    defparam I1.init = 16'b0000000011111111;
    
endmodule
//
// Verilog Description of module inverter_U57
//

module inverter_U57 (\notGate[947]_keep , \notGate[948] ) /* synthesis syn_module_defined=1 */ ;
    input \notGate[947]_keep ;
    output \notGate[948] ;
    
    wire \notGate[947]_keep  /* synthesis alspreserve=1 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(25[15:22])
    
    LUT4 I1 (.A(\notGate[947]_keep ), .B(\notGate[947]_keep ), .C(\notGate[947]_keep ), 
         .D(\notGate[947]_keep ), .Z(\notGate[948] )) /* synthesis syn_instantiated=1, lut_function=((!D !C !B !A)+(!D !C !B A)+(!D !C B !A)+(!D !C B A)+(!D C !B !A)+(!D C !B A)+(!D C B !A)+(!D C B A)), LSE_LINE_FILE_ID=3, LSE_LCOL=13, LSE_RCOL=44, LSE_LLINE=32, LSE_RLINE=32 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(11[2:53])
    defparam I1.init = 16'b0000000011111111;
    
endmodule
//
// Verilog Description of module inverter_U58
//

module inverter_U58 (\notGate[946]_keep , \notGate[947] ) /* synthesis syn_module_defined=1 */ ;
    input \notGate[946]_keep ;
    output \notGate[947] ;
    
    wire \notGate[946]_keep  /* synthesis alspreserve=1 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(25[15:22])
    
    LUT4 I1 (.A(\notGate[946]_keep ), .B(\notGate[946]_keep ), .C(\notGate[946]_keep ), 
         .D(\notGate[946]_keep ), .Z(\notGate[947] )) /* synthesis syn_instantiated=1, lut_function=((!D !C !B !A)+(!D !C !B A)+(!D !C B !A)+(!D !C B A)+(!D C !B !A)+(!D C !B A)+(!D C B !A)+(!D C B A)), LSE_LINE_FILE_ID=3, LSE_LCOL=13, LSE_RCOL=44, LSE_LLINE=32, LSE_RLINE=32 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(11[2:53])
    defparam I1.init = 16'b0000000011111111;
    
endmodule
//
// Verilog Description of module inverter_U59
//

module inverter_U59 (\notGate[945]_keep , \notGate[946] ) /* synthesis syn_module_defined=1 */ ;
    input \notGate[945]_keep ;
    output \notGate[946] ;
    
    wire \notGate[945]_keep  /* synthesis alspreserve=1 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(25[15:22])
    
    LUT4 I1 (.A(\notGate[945]_keep ), .B(\notGate[945]_keep ), .C(\notGate[945]_keep ), 
         .D(\notGate[945]_keep ), .Z(\notGate[946] )) /* synthesis syn_instantiated=1, lut_function=((!D !C !B !A)+(!D !C !B A)+(!D !C B !A)+(!D !C B A)+(!D C !B !A)+(!D C !B A)+(!D C B !A)+(!D C B A)), LSE_LINE_FILE_ID=3, LSE_LCOL=13, LSE_RCOL=44, LSE_LLINE=32, LSE_RLINE=32 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(11[2:53])
    defparam I1.init = 16'b0000000011111111;
    
endmodule
//
// Verilog Description of module inverter_U60
//

module inverter_U60 (\notGate[944]_keep , \notGate[945] ) /* synthesis syn_module_defined=1 */ ;
    input \notGate[944]_keep ;
    output \notGate[945] ;
    
    wire \notGate[944]_keep  /* synthesis alspreserve=1 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(25[15:22])
    
    LUT4 I1 (.A(\notGate[944]_keep ), .B(\notGate[944]_keep ), .C(\notGate[944]_keep ), 
         .D(\notGate[944]_keep ), .Z(\notGate[945] )) /* synthesis syn_instantiated=1, lut_function=((!D !C !B !A)+(!D !C !B A)+(!D !C B !A)+(!D !C B A)+(!D C !B !A)+(!D C !B A)+(!D C B !A)+(!D C B A)), LSE_LINE_FILE_ID=3, LSE_LCOL=13, LSE_RCOL=44, LSE_LLINE=32, LSE_RLINE=32 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(11[2:53])
    defparam I1.init = 16'b0000000011111111;
    
endmodule
//
// Verilog Description of module inverter_U61
//

module inverter_U61 (\notGate[943]_keep , \notGate[944] ) /* synthesis syn_module_defined=1 */ ;
    input \notGate[943]_keep ;
    output \notGate[944] ;
    
    wire \notGate[943]_keep  /* synthesis alspreserve=1 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(25[15:22])
    
    LUT4 I1 (.A(\notGate[943]_keep ), .B(\notGate[943]_keep ), .C(\notGate[943]_keep ), 
         .D(\notGate[943]_keep ), .Z(\notGate[944] )) /* synthesis syn_instantiated=1, lut_function=((!D !C !B !A)+(!D !C !B A)+(!D !C B !A)+(!D !C B A)+(!D C !B !A)+(!D C !B A)+(!D C B !A)+(!D C B A)), LSE_LINE_FILE_ID=3, LSE_LCOL=13, LSE_RCOL=44, LSE_LLINE=32, LSE_RLINE=32 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(11[2:53])
    defparam I1.init = 16'b0000000011111111;
    
endmodule
//
// Verilog Description of module inverter_U62
//

module inverter_U62 (\notGate[942]_keep , \notGate[943] ) /* synthesis syn_module_defined=1 */ ;
    input \notGate[942]_keep ;
    output \notGate[943] ;
    
    wire \notGate[942]_keep  /* synthesis alspreserve=1 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(25[15:22])
    
    LUT4 I1 (.A(\notGate[942]_keep ), .B(\notGate[942]_keep ), .C(\notGate[942]_keep ), 
         .D(\notGate[942]_keep ), .Z(\notGate[943] )) /* synthesis syn_instantiated=1, lut_function=((!D !C !B !A)+(!D !C !B A)+(!D !C B !A)+(!D !C B A)+(!D C !B !A)+(!D C !B A)+(!D C B !A)+(!D C B A)), LSE_LINE_FILE_ID=3, LSE_LCOL=13, LSE_RCOL=44, LSE_LLINE=32, LSE_RLINE=32 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(11[2:53])
    defparam I1.init = 16'b0000000011111111;
    
endmodule
//
// Verilog Description of module inverter_U63
//

module inverter_U63 (\notGate[941]_keep , \notGate[942] ) /* synthesis syn_module_defined=1 */ ;
    input \notGate[941]_keep ;
    output \notGate[942] ;
    
    wire \notGate[941]_keep  /* synthesis alspreserve=1 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(25[15:22])
    
    LUT4 I1 (.A(\notGate[941]_keep ), .B(\notGate[941]_keep ), .C(\notGate[941]_keep ), 
         .D(\notGate[941]_keep ), .Z(\notGate[942] )) /* synthesis syn_instantiated=1, lut_function=((!D !C !B !A)+(!D !C !B A)+(!D !C B !A)+(!D !C B A)+(!D C !B !A)+(!D C !B A)+(!D C B !A)+(!D C B A)), LSE_LINE_FILE_ID=3, LSE_LCOL=13, LSE_RCOL=44, LSE_LLINE=32, LSE_RLINE=32 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(11[2:53])
    defparam I1.init = 16'b0000000011111111;
    
endmodule
//
// Verilog Description of module inverter_U64
//

module inverter_U64 (\notGate[940]_keep , \notGate[941] ) /* synthesis syn_module_defined=1 */ ;
    input \notGate[940]_keep ;
    output \notGate[941] ;
    
    wire \notGate[940]_keep  /* synthesis alspreserve=1 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(25[15:22])
    
    LUT4 I1 (.A(\notGate[940]_keep ), .B(\notGate[940]_keep ), .C(\notGate[940]_keep ), 
         .D(\notGate[940]_keep ), .Z(\notGate[941] )) /* synthesis syn_instantiated=1, lut_function=((!D !C !B !A)+(!D !C !B A)+(!D !C B !A)+(!D !C B A)+(!D C !B !A)+(!D C !B A)+(!D C B !A)+(!D C B A)), LSE_LINE_FILE_ID=3, LSE_LCOL=13, LSE_RCOL=44, LSE_LLINE=32, LSE_RLINE=32 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(11[2:53])
    defparam I1.init = 16'b0000000011111111;
    
endmodule
//
// Verilog Description of module inverter_U65
//

module inverter_U65 (\notGate[939]_keep , \notGate[940] ) /* synthesis syn_module_defined=1 */ ;
    input \notGate[939]_keep ;
    output \notGate[940] ;
    
    wire \notGate[939]_keep  /* synthesis alspreserve=1 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(25[15:22])
    
    LUT4 I1 (.A(\notGate[939]_keep ), .B(\notGate[939]_keep ), .C(\notGate[939]_keep ), 
         .D(\notGate[939]_keep ), .Z(\notGate[940] )) /* synthesis syn_instantiated=1, lut_function=((!D !C !B !A)+(!D !C !B A)+(!D !C B !A)+(!D !C B A)+(!D C !B !A)+(!D C !B A)+(!D C B !A)+(!D C B A)), LSE_LINE_FILE_ID=3, LSE_LCOL=13, LSE_RCOL=44, LSE_LLINE=32, LSE_RLINE=32 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(11[2:53])
    defparam I1.init = 16'b0000000011111111;
    
endmodule
//
// Verilog Description of module inverter_U66
//

module inverter_U66 (\notGate[92]_keep , \notGate[93] ) /* synthesis syn_module_defined=1 */ ;
    input \notGate[92]_keep ;
    output \notGate[93] ;
    
    wire \notGate[92]_keep  /* synthesis alspreserve=1 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(25[15:22])
    
    LUT4 I1 (.A(\notGate[92]_keep ), .B(\notGate[92]_keep ), .C(\notGate[92]_keep ), 
         .D(\notGate[92]_keep ), .Z(\notGate[93] )) /* synthesis syn_instantiated=1, lut_function=((!D !C !B !A)+(!D !C !B A)+(!D !C B !A)+(!D !C B A)+(!D C !B !A)+(!D C !B A)+(!D C B !A)+(!D C B A)), LSE_LINE_FILE_ID=3, LSE_LCOL=13, LSE_RCOL=44, LSE_LLINE=32, LSE_RLINE=32 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(11[2:53])
    defparam I1.init = 16'b0000000011111111;
    
endmodule
//
// Verilog Description of module inverter_U67
//

module inverter_U67 (\notGate[938]_keep , \notGate[939] ) /* synthesis syn_module_defined=1 */ ;
    input \notGate[938]_keep ;
    output \notGate[939] ;
    
    wire \notGate[938]_keep  /* synthesis alspreserve=1 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(25[15:22])
    
    LUT4 I1 (.A(\notGate[938]_keep ), .B(\notGate[938]_keep ), .C(\notGate[938]_keep ), 
         .D(\notGate[938]_keep ), .Z(\notGate[939] )) /* synthesis syn_instantiated=1, lut_function=((!D !C !B !A)+(!D !C !B A)+(!D !C B !A)+(!D !C B A)+(!D C !B !A)+(!D C !B A)+(!D C B !A)+(!D C B A)), LSE_LINE_FILE_ID=3, LSE_LCOL=13, LSE_RCOL=44, LSE_LLINE=32, LSE_RLINE=32 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(11[2:53])
    defparam I1.init = 16'b0000000011111111;
    
endmodule
//
// Verilog Description of module inverter_U68
//

module inverter_U68 (\notGate[937]_keep , \notGate[938] ) /* synthesis syn_module_defined=1 */ ;
    input \notGate[937]_keep ;
    output \notGate[938] ;
    
    wire \notGate[937]_keep  /* synthesis alspreserve=1 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(25[15:22])
    
    LUT4 I1 (.A(\notGate[937]_keep ), .B(\notGate[937]_keep ), .C(\notGate[937]_keep ), 
         .D(\notGate[937]_keep ), .Z(\notGate[938] )) /* synthesis syn_instantiated=1, lut_function=((!D !C !B !A)+(!D !C !B A)+(!D !C B !A)+(!D !C B A)+(!D C !B !A)+(!D C !B A)+(!D C B !A)+(!D C B A)), LSE_LINE_FILE_ID=3, LSE_LCOL=13, LSE_RCOL=44, LSE_LLINE=32, LSE_RLINE=32 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(11[2:53])
    defparam I1.init = 16'b0000000011111111;
    
endmodule
//
// Verilog Description of module inverter_U69
//

module inverter_U69 (\notGate[936]_keep , \notGate[937] ) /* synthesis syn_module_defined=1 */ ;
    input \notGate[936]_keep ;
    output \notGate[937] ;
    
    wire \notGate[936]_keep  /* synthesis alspreserve=1 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(25[15:22])
    
    LUT4 I1 (.A(\notGate[936]_keep ), .B(\notGate[936]_keep ), .C(\notGate[936]_keep ), 
         .D(\notGate[936]_keep ), .Z(\notGate[937] )) /* synthesis syn_instantiated=1, lut_function=((!D !C !B !A)+(!D !C !B A)+(!D !C B !A)+(!D !C B A)+(!D C !B !A)+(!D C !B A)+(!D C B !A)+(!D C B A)), LSE_LINE_FILE_ID=3, LSE_LCOL=13, LSE_RCOL=44, LSE_LLINE=32, LSE_RLINE=32 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(11[2:53])
    defparam I1.init = 16'b0000000011111111;
    
endmodule
//
// Verilog Description of module inverter_U70
//

module inverter_U70 (\notGate[935]_keep , \notGate[936] ) /* synthesis syn_module_defined=1 */ ;
    input \notGate[935]_keep ;
    output \notGate[936] ;
    
    wire \notGate[935]_keep  /* synthesis alspreserve=1 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(25[15:22])
    
    LUT4 I1 (.A(\notGate[935]_keep ), .B(\notGate[935]_keep ), .C(\notGate[935]_keep ), 
         .D(\notGate[935]_keep ), .Z(\notGate[936] )) /* synthesis syn_instantiated=1, lut_function=((!D !C !B !A)+(!D !C !B A)+(!D !C B !A)+(!D !C B A)+(!D C !B !A)+(!D C !B A)+(!D C B !A)+(!D C B A)), LSE_LINE_FILE_ID=3, LSE_LCOL=13, LSE_RCOL=44, LSE_LLINE=32, LSE_RLINE=32 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(11[2:53])
    defparam I1.init = 16'b0000000011111111;
    
endmodule
//
// Verilog Description of module inverter_U71
//

module inverter_U71 (\notGate[934]_keep , \notGate[935] ) /* synthesis syn_module_defined=1 */ ;
    input \notGate[934]_keep ;
    output \notGate[935] ;
    
    wire \notGate[934]_keep  /* synthesis alspreserve=1 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(25[15:22])
    
    LUT4 I1 (.A(\notGate[934]_keep ), .B(\notGate[934]_keep ), .C(\notGate[934]_keep ), 
         .D(\notGate[934]_keep ), .Z(\notGate[935] )) /* synthesis syn_instantiated=1, lut_function=((!D !C !B !A)+(!D !C !B A)+(!D !C B !A)+(!D !C B A)+(!D C !B !A)+(!D C !B A)+(!D C B !A)+(!D C B A)), LSE_LINE_FILE_ID=3, LSE_LCOL=13, LSE_RCOL=44, LSE_LLINE=32, LSE_RLINE=32 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(11[2:53])
    defparam I1.init = 16'b0000000011111111;
    
endmodule
//
// Verilog Description of module inverter_U72
//

module inverter_U72 (\notGate[933]_keep , \notGate[934] ) /* synthesis syn_module_defined=1 */ ;
    input \notGate[933]_keep ;
    output \notGate[934] ;
    
    wire \notGate[933]_keep  /* synthesis alspreserve=1 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(25[15:22])
    
    LUT4 I1 (.A(\notGate[933]_keep ), .B(\notGate[933]_keep ), .C(\notGate[933]_keep ), 
         .D(\notGate[933]_keep ), .Z(\notGate[934] )) /* synthesis syn_instantiated=1, lut_function=((!D !C !B !A)+(!D !C !B A)+(!D !C B !A)+(!D !C B A)+(!D C !B !A)+(!D C !B A)+(!D C B !A)+(!D C B A)), LSE_LINE_FILE_ID=3, LSE_LCOL=13, LSE_RCOL=44, LSE_LLINE=32, LSE_RLINE=32 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(11[2:53])
    defparam I1.init = 16'b0000000011111111;
    
endmodule
//
// Verilog Description of module inverter_U73
//

module inverter_U73 (\notGate[932]_keep , \notGate[933] ) /* synthesis syn_module_defined=1 */ ;
    input \notGate[932]_keep ;
    output \notGate[933] ;
    
    wire \notGate[932]_keep  /* synthesis alspreserve=1 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(25[15:22])
    
    LUT4 I1 (.A(\notGate[932]_keep ), .B(\notGate[932]_keep ), .C(\notGate[932]_keep ), 
         .D(\notGate[932]_keep ), .Z(\notGate[933] )) /* synthesis syn_instantiated=1, lut_function=((!D !C !B !A)+(!D !C !B A)+(!D !C B !A)+(!D !C B A)+(!D C !B !A)+(!D C !B A)+(!D C B !A)+(!D C B A)), LSE_LINE_FILE_ID=3, LSE_LCOL=13, LSE_RCOL=44, LSE_LLINE=32, LSE_RLINE=32 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(11[2:53])
    defparam I1.init = 16'b0000000011111111;
    
endmodule
//
// Verilog Description of module inverter_U74
//

module inverter_U74 (\notGate[931]_keep , \notGate[932] ) /* synthesis syn_module_defined=1 */ ;
    input \notGate[931]_keep ;
    output \notGate[932] ;
    
    wire \notGate[931]_keep  /* synthesis alspreserve=1 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(25[15:22])
    
    LUT4 I1 (.A(\notGate[931]_keep ), .B(\notGate[931]_keep ), .C(\notGate[931]_keep ), 
         .D(\notGate[931]_keep ), .Z(\notGate[932] )) /* synthesis syn_instantiated=1, lut_function=((!D !C !B !A)+(!D !C !B A)+(!D !C B !A)+(!D !C B A)+(!D C !B !A)+(!D C !B A)+(!D C B !A)+(!D C B A)), LSE_LINE_FILE_ID=3, LSE_LCOL=13, LSE_RCOL=44, LSE_LLINE=32, LSE_RLINE=32 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(11[2:53])
    defparam I1.init = 16'b0000000011111111;
    
endmodule
//
// Verilog Description of module inverter_U75
//

module inverter_U75 (\notGate[930]_keep , \notGate[931] ) /* synthesis syn_module_defined=1 */ ;
    input \notGate[930]_keep ;
    output \notGate[931] ;
    
    wire \notGate[930]_keep  /* synthesis alspreserve=1 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(25[15:22])
    
    LUT4 I1 (.A(\notGate[930]_keep ), .B(\notGate[930]_keep ), .C(\notGate[930]_keep ), 
         .D(\notGate[930]_keep ), .Z(\notGate[931] )) /* synthesis syn_instantiated=1, lut_function=((!D !C !B !A)+(!D !C !B A)+(!D !C B !A)+(!D !C B A)+(!D C !B !A)+(!D C !B A)+(!D C B !A)+(!D C B A)), LSE_LINE_FILE_ID=3, LSE_LCOL=13, LSE_RCOL=44, LSE_LLINE=32, LSE_RLINE=32 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(11[2:53])
    defparam I1.init = 16'b0000000011111111;
    
endmodule
//
// Verilog Description of module inverter_U76
//

module inverter_U76 (\notGate[929]_keep , \notGate[930] ) /* synthesis syn_module_defined=1 */ ;
    input \notGate[929]_keep ;
    output \notGate[930] ;
    
    wire \notGate[929]_keep  /* synthesis alspreserve=1 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(25[15:22])
    
    LUT4 I1 (.A(\notGate[929]_keep ), .B(\notGate[929]_keep ), .C(\notGate[929]_keep ), 
         .D(\notGate[929]_keep ), .Z(\notGate[930] )) /* synthesis syn_instantiated=1, lut_function=((!D !C !B !A)+(!D !C !B A)+(!D !C B !A)+(!D !C B A)+(!D C !B !A)+(!D C !B A)+(!D C B !A)+(!D C B A)), LSE_LINE_FILE_ID=3, LSE_LCOL=13, LSE_RCOL=44, LSE_LLINE=32, LSE_RLINE=32 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(11[2:53])
    defparam I1.init = 16'b0000000011111111;
    
endmodule
//
// Verilog Description of module inverter_U77
//

module inverter_U77 (\notGate[91]_keep , \notGate[92] ) /* synthesis syn_module_defined=1 */ ;
    input \notGate[91]_keep ;
    output \notGate[92] ;
    
    wire \notGate[91]_keep  /* synthesis alspreserve=1 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(25[15:22])
    
    LUT4 I1 (.A(\notGate[91]_keep ), .B(\notGate[91]_keep ), .C(\notGate[91]_keep ), 
         .D(\notGate[91]_keep ), .Z(\notGate[92] )) /* synthesis syn_instantiated=1, lut_function=((!D !C !B !A)+(!D !C !B A)+(!D !C B !A)+(!D !C B A)+(!D C !B !A)+(!D C !B A)+(!D C B !A)+(!D C B A)), LSE_LINE_FILE_ID=3, LSE_LCOL=13, LSE_RCOL=44, LSE_LLINE=32, LSE_RLINE=32 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(11[2:53])
    defparam I1.init = 16'b0000000011111111;
    
endmodule
//
// Verilog Description of module inverter_U78
//

module inverter_U78 (\notGate[928]_keep , \notGate[929] ) /* synthesis syn_module_defined=1 */ ;
    input \notGate[928]_keep ;
    output \notGate[929] ;
    
    wire \notGate[928]_keep  /* synthesis alspreserve=1 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(25[15:22])
    
    LUT4 I1 (.A(\notGate[928]_keep ), .B(\notGate[928]_keep ), .C(\notGate[928]_keep ), 
         .D(\notGate[928]_keep ), .Z(\notGate[929] )) /* synthesis syn_instantiated=1, lut_function=((!D !C !B !A)+(!D !C !B A)+(!D !C B !A)+(!D !C B A)+(!D C !B !A)+(!D C !B A)+(!D C B !A)+(!D C B A)), LSE_LINE_FILE_ID=3, LSE_LCOL=13, LSE_RCOL=44, LSE_LLINE=32, LSE_RLINE=32 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(11[2:53])
    defparam I1.init = 16'b0000000011111111;
    
endmodule
//
// Verilog Description of module inverter_U79
//

module inverter_U79 (\notGate[927]_keep , \notGate[928] ) /* synthesis syn_module_defined=1 */ ;
    input \notGate[927]_keep ;
    output \notGate[928] ;
    
    wire \notGate[927]_keep  /* synthesis alspreserve=1 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(25[15:22])
    
    LUT4 I1 (.A(\notGate[927]_keep ), .B(\notGate[927]_keep ), .C(\notGate[927]_keep ), 
         .D(\notGate[927]_keep ), .Z(\notGate[928] )) /* synthesis syn_instantiated=1, lut_function=((!D !C !B !A)+(!D !C !B A)+(!D !C B !A)+(!D !C B A)+(!D C !B !A)+(!D C !B A)+(!D C B !A)+(!D C B A)), LSE_LINE_FILE_ID=3, LSE_LCOL=13, LSE_RCOL=44, LSE_LLINE=32, LSE_RLINE=32 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(11[2:53])
    defparam I1.init = 16'b0000000011111111;
    
endmodule
//
// Verilog Description of module inverter_U80
//

module inverter_U80 (\notGate[926]_keep , \notGate[927] ) /* synthesis syn_module_defined=1 */ ;
    input \notGate[926]_keep ;
    output \notGate[927] ;
    
    wire \notGate[926]_keep  /* synthesis alspreserve=1 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(25[15:22])
    
    LUT4 I1 (.A(\notGate[926]_keep ), .B(\notGate[926]_keep ), .C(\notGate[926]_keep ), 
         .D(\notGate[926]_keep ), .Z(\notGate[927] )) /* synthesis syn_instantiated=1, lut_function=((!D !C !B !A)+(!D !C !B A)+(!D !C B !A)+(!D !C B A)+(!D C !B !A)+(!D C !B A)+(!D C B !A)+(!D C B A)), LSE_LINE_FILE_ID=3, LSE_LCOL=13, LSE_RCOL=44, LSE_LLINE=32, LSE_RLINE=32 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(11[2:53])
    defparam I1.init = 16'b0000000011111111;
    
endmodule
//
// Verilog Description of module inverter_U81
//

module inverter_U81 (\notGate[925]_keep , \notGate[926] ) /* synthesis syn_module_defined=1 */ ;
    input \notGate[925]_keep ;
    output \notGate[926] ;
    
    wire \notGate[925]_keep  /* synthesis alspreserve=1 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(25[15:22])
    
    LUT4 I1 (.A(\notGate[925]_keep ), .B(\notGate[925]_keep ), .C(\notGate[925]_keep ), 
         .D(\notGate[925]_keep ), .Z(\notGate[926] )) /* synthesis syn_instantiated=1, lut_function=((!D !C !B !A)+(!D !C !B A)+(!D !C B !A)+(!D !C B A)+(!D C !B !A)+(!D C !B A)+(!D C B !A)+(!D C B A)), LSE_LINE_FILE_ID=3, LSE_LCOL=13, LSE_RCOL=44, LSE_LLINE=32, LSE_RLINE=32 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(11[2:53])
    defparam I1.init = 16'b0000000011111111;
    
endmodule
//
// Verilog Description of module inverter_U82
//

module inverter_U82 (\notGate[924]_keep , \notGate[925] ) /* synthesis syn_module_defined=1 */ ;
    input \notGate[924]_keep ;
    output \notGate[925] ;
    
    wire \notGate[924]_keep  /* synthesis alspreserve=1 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(25[15:22])
    
    LUT4 I1 (.A(\notGate[924]_keep ), .B(\notGate[924]_keep ), .C(\notGate[924]_keep ), 
         .D(\notGate[924]_keep ), .Z(\notGate[925] )) /* synthesis syn_instantiated=1, lut_function=((!D !C !B !A)+(!D !C !B A)+(!D !C B !A)+(!D !C B A)+(!D C !B !A)+(!D C !B A)+(!D C B !A)+(!D C B A)), LSE_LINE_FILE_ID=3, LSE_LCOL=13, LSE_RCOL=44, LSE_LLINE=32, LSE_RLINE=32 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(11[2:53])
    defparam I1.init = 16'b0000000011111111;
    
endmodule
//
// Verilog Description of module inverter_U83
//

module inverter_U83 (\notGate[923]_keep , \notGate[924] ) /* synthesis syn_module_defined=1 */ ;
    input \notGate[923]_keep ;
    output \notGate[924] ;
    
    wire \notGate[923]_keep  /* synthesis alspreserve=1 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(25[15:22])
    
    LUT4 I1 (.A(\notGate[923]_keep ), .B(\notGate[923]_keep ), .C(\notGate[923]_keep ), 
         .D(\notGate[923]_keep ), .Z(\notGate[924] )) /* synthesis syn_instantiated=1, lut_function=((!D !C !B !A)+(!D !C !B A)+(!D !C B !A)+(!D !C B A)+(!D C !B !A)+(!D C !B A)+(!D C B !A)+(!D C B A)), LSE_LINE_FILE_ID=3, LSE_LCOL=13, LSE_RCOL=44, LSE_LLINE=32, LSE_RLINE=32 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(11[2:53])
    defparam I1.init = 16'b0000000011111111;
    
endmodule
//
// Verilog Description of module inverter_U84
//

module inverter_U84 (\notGate[922]_keep , \notGate[923] ) /* synthesis syn_module_defined=1 */ ;
    input \notGate[922]_keep ;
    output \notGate[923] ;
    
    wire \notGate[922]_keep  /* synthesis alspreserve=1 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(25[15:22])
    
    LUT4 I1 (.A(\notGate[922]_keep ), .B(\notGate[922]_keep ), .C(\notGate[922]_keep ), 
         .D(\notGate[922]_keep ), .Z(\notGate[923] )) /* synthesis syn_instantiated=1, lut_function=((!D !C !B !A)+(!D !C !B A)+(!D !C B !A)+(!D !C B A)+(!D C !B !A)+(!D C !B A)+(!D C B !A)+(!D C B A)), LSE_LINE_FILE_ID=3, LSE_LCOL=13, LSE_RCOL=44, LSE_LLINE=32, LSE_RLINE=32 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(11[2:53])
    defparam I1.init = 16'b0000000011111111;
    
endmodule
//
// Verilog Description of module inverter_U85
//

module inverter_U85 (\notGate[921]_keep , \notGate[922] ) /* synthesis syn_module_defined=1 */ ;
    input \notGate[921]_keep ;
    output \notGate[922] ;
    
    wire \notGate[921]_keep  /* synthesis alspreserve=1 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(25[15:22])
    
    LUT4 I1 (.A(\notGate[921]_keep ), .B(\notGate[921]_keep ), .C(\notGate[921]_keep ), 
         .D(\notGate[921]_keep ), .Z(\notGate[922] )) /* synthesis syn_instantiated=1, lut_function=((!D !C !B !A)+(!D !C !B A)+(!D !C B !A)+(!D !C B A)+(!D C !B !A)+(!D C !B A)+(!D C B !A)+(!D C B A)), LSE_LINE_FILE_ID=3, LSE_LCOL=13, LSE_RCOL=44, LSE_LLINE=32, LSE_RLINE=32 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(11[2:53])
    defparam I1.init = 16'b0000000011111111;
    
endmodule
//
// Verilog Description of module inverter_U86
//

module inverter_U86 (\notGate[920]_keep , \notGate[921] ) /* synthesis syn_module_defined=1 */ ;
    input \notGate[920]_keep ;
    output \notGate[921] ;
    
    wire \notGate[920]_keep  /* synthesis alspreserve=1 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(25[15:22])
    
    LUT4 I1 (.A(\notGate[920]_keep ), .B(\notGate[920]_keep ), .C(\notGate[920]_keep ), 
         .D(\notGate[920]_keep ), .Z(\notGate[921] )) /* synthesis syn_instantiated=1, lut_function=((!D !C !B !A)+(!D !C !B A)+(!D !C B !A)+(!D !C B A)+(!D C !B !A)+(!D C !B A)+(!D C B !A)+(!D C B A)), LSE_LINE_FILE_ID=3, LSE_LCOL=13, LSE_RCOL=44, LSE_LLINE=32, LSE_RLINE=32 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(11[2:53])
    defparam I1.init = 16'b0000000011111111;
    
endmodule
//
// Verilog Description of module inverter_U87
//

module inverter_U87 (\notGate[919]_keep , \notGate[920] ) /* synthesis syn_module_defined=1 */ ;
    input \notGate[919]_keep ;
    output \notGate[920] ;
    
    wire \notGate[919]_keep  /* synthesis alspreserve=1 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(25[15:22])
    
    LUT4 I1 (.A(\notGate[919]_keep ), .B(\notGate[919]_keep ), .C(\notGate[919]_keep ), 
         .D(\notGate[919]_keep ), .Z(\notGate[920] )) /* synthesis syn_instantiated=1, lut_function=((!D !C !B !A)+(!D !C !B A)+(!D !C B !A)+(!D !C B A)+(!D C !B !A)+(!D C !B A)+(!D C B !A)+(!D C B A)), LSE_LINE_FILE_ID=3, LSE_LCOL=13, LSE_RCOL=44, LSE_LLINE=32, LSE_RLINE=32 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(11[2:53])
    defparam I1.init = 16'b0000000011111111;
    
endmodule
//
// Verilog Description of module inverter_U88
//

module inverter_U88 (\notGate[90]_keep , \notGate[91] ) /* synthesis syn_module_defined=1 */ ;
    input \notGate[90]_keep ;
    output \notGate[91] ;
    
    wire \notGate[90]_keep  /* synthesis alspreserve=1 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(25[15:22])
    
    LUT4 I1 (.A(\notGate[90]_keep ), .B(\notGate[90]_keep ), .C(\notGate[90]_keep ), 
         .D(\notGate[90]_keep ), .Z(\notGate[91] )) /* synthesis syn_instantiated=1, lut_function=((!D !C !B !A)+(!D !C !B A)+(!D !C B !A)+(!D !C B A)+(!D C !B !A)+(!D C !B A)+(!D C B !A)+(!D C B A)), LSE_LINE_FILE_ID=3, LSE_LCOL=13, LSE_RCOL=44, LSE_LLINE=32, LSE_RLINE=32 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(11[2:53])
    defparam I1.init = 16'b0000000011111111;
    
endmodule
//
// Verilog Description of module inverter_U89
//

module inverter_U89 (\notGate[918]_keep , \notGate[919] ) /* synthesis syn_module_defined=1 */ ;
    input \notGate[918]_keep ;
    output \notGate[919] ;
    
    wire \notGate[918]_keep  /* synthesis alspreserve=1 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(25[15:22])
    
    LUT4 I1 (.A(\notGate[918]_keep ), .B(\notGate[918]_keep ), .C(\notGate[918]_keep ), 
         .D(\notGate[918]_keep ), .Z(\notGate[919] )) /* synthesis syn_instantiated=1, lut_function=((!D !C !B !A)+(!D !C !B A)+(!D !C B !A)+(!D !C B A)+(!D C !B !A)+(!D C !B A)+(!D C B !A)+(!D C B A)), LSE_LINE_FILE_ID=3, LSE_LCOL=13, LSE_RCOL=44, LSE_LLINE=32, LSE_RLINE=32 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(11[2:53])
    defparam I1.init = 16'b0000000011111111;
    
endmodule
//
// Verilog Description of module inverter_U90
//

module inverter_U90 (\notGate[917]_keep , \notGate[918] ) /* synthesis syn_module_defined=1 */ ;
    input \notGate[917]_keep ;
    output \notGate[918] ;
    
    wire \notGate[917]_keep  /* synthesis alspreserve=1 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(25[15:22])
    
    LUT4 I1 (.A(\notGate[917]_keep ), .B(\notGate[917]_keep ), .C(\notGate[917]_keep ), 
         .D(\notGate[917]_keep ), .Z(\notGate[918] )) /* synthesis syn_instantiated=1, lut_function=((!D !C !B !A)+(!D !C !B A)+(!D !C B !A)+(!D !C B A)+(!D C !B !A)+(!D C !B A)+(!D C B !A)+(!D C B A)), LSE_LINE_FILE_ID=3, LSE_LCOL=13, LSE_RCOL=44, LSE_LLINE=32, LSE_RLINE=32 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(11[2:53])
    defparam I1.init = 16'b0000000011111111;
    
endmodule
//
// Verilog Description of module inverter_U91
//

module inverter_U91 (\notGate[916]_keep , \notGate[917] ) /* synthesis syn_module_defined=1 */ ;
    input \notGate[916]_keep ;
    output \notGate[917] ;
    
    wire \notGate[916]_keep  /* synthesis alspreserve=1 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(25[15:22])
    
    LUT4 I1 (.A(\notGate[916]_keep ), .B(\notGate[916]_keep ), .C(\notGate[916]_keep ), 
         .D(\notGate[916]_keep ), .Z(\notGate[917] )) /* synthesis syn_instantiated=1, lut_function=((!D !C !B !A)+(!D !C !B A)+(!D !C B !A)+(!D !C B A)+(!D C !B !A)+(!D C !B A)+(!D C B !A)+(!D C B A)), LSE_LINE_FILE_ID=3, LSE_LCOL=13, LSE_RCOL=44, LSE_LLINE=32, LSE_RLINE=32 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(11[2:53])
    defparam I1.init = 16'b0000000011111111;
    
endmodule
//
// Verilog Description of module inverter_U92
//

module inverter_U92 (\notGate[915]_keep , \notGate[916] ) /* synthesis syn_module_defined=1 */ ;
    input \notGate[915]_keep ;
    output \notGate[916] ;
    
    wire \notGate[915]_keep  /* synthesis alspreserve=1 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(25[15:22])
    
    LUT4 I1 (.A(\notGate[915]_keep ), .B(\notGate[915]_keep ), .C(\notGate[915]_keep ), 
         .D(\notGate[915]_keep ), .Z(\notGate[916] )) /* synthesis syn_instantiated=1, lut_function=((!D !C !B !A)+(!D !C !B A)+(!D !C B !A)+(!D !C B A)+(!D C !B !A)+(!D C !B A)+(!D C B !A)+(!D C B A)), LSE_LINE_FILE_ID=3, LSE_LCOL=13, LSE_RCOL=44, LSE_LLINE=32, LSE_RLINE=32 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(11[2:53])
    defparam I1.init = 16'b0000000011111111;
    
endmodule
//
// Verilog Description of module inverter_U93
//

module inverter_U93 (\notGate[914]_keep , \notGate[915] ) /* synthesis syn_module_defined=1 */ ;
    input \notGate[914]_keep ;
    output \notGate[915] ;
    
    wire \notGate[914]_keep  /* synthesis alspreserve=1 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(25[15:22])
    
    LUT4 I1 (.A(\notGate[914]_keep ), .B(\notGate[914]_keep ), .C(\notGate[914]_keep ), 
         .D(\notGate[914]_keep ), .Z(\notGate[915] )) /* synthesis syn_instantiated=1, lut_function=((!D !C !B !A)+(!D !C !B A)+(!D !C B !A)+(!D !C B A)+(!D C !B !A)+(!D C !B A)+(!D C B !A)+(!D C B A)), LSE_LINE_FILE_ID=3, LSE_LCOL=13, LSE_RCOL=44, LSE_LLINE=32, LSE_RLINE=32 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(11[2:53])
    defparam I1.init = 16'b0000000011111111;
    
endmodule
//
// Verilog Description of module inverter_U94
//

module inverter_U94 (\notGate[913]_keep , \notGate[914] ) /* synthesis syn_module_defined=1 */ ;
    input \notGate[913]_keep ;
    output \notGate[914] ;
    
    wire \notGate[913]_keep  /* synthesis alspreserve=1 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(25[15:22])
    
    LUT4 I1 (.A(\notGate[913]_keep ), .B(\notGate[913]_keep ), .C(\notGate[913]_keep ), 
         .D(\notGate[913]_keep ), .Z(\notGate[914] )) /* synthesis syn_instantiated=1, lut_function=((!D !C !B !A)+(!D !C !B A)+(!D !C B !A)+(!D !C B A)+(!D C !B !A)+(!D C !B A)+(!D C B !A)+(!D C B A)), LSE_LINE_FILE_ID=3, LSE_LCOL=13, LSE_RCOL=44, LSE_LLINE=32, LSE_RLINE=32 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(11[2:53])
    defparam I1.init = 16'b0000000011111111;
    
endmodule
//
// Verilog Description of module inverter_U95
//

module inverter_U95 (\notGate[912]_keep , \notGate[913] ) /* synthesis syn_module_defined=1 */ ;
    input \notGate[912]_keep ;
    output \notGate[913] ;
    
    wire \notGate[912]_keep  /* synthesis alspreserve=1 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(25[15:22])
    
    LUT4 I1 (.A(\notGate[912]_keep ), .B(\notGate[912]_keep ), .C(\notGate[912]_keep ), 
         .D(\notGate[912]_keep ), .Z(\notGate[913] )) /* synthesis syn_instantiated=1, lut_function=((!D !C !B !A)+(!D !C !B A)+(!D !C B !A)+(!D !C B A)+(!D C !B !A)+(!D C !B A)+(!D C B !A)+(!D C B A)), LSE_LINE_FILE_ID=3, LSE_LCOL=13, LSE_RCOL=44, LSE_LLINE=32, LSE_RLINE=32 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(11[2:53])
    defparam I1.init = 16'b0000000011111111;
    
endmodule
//
// Verilog Description of module inverter_U96
//

module inverter_U96 (\notGate[911]_keep , \notGate[912] ) /* synthesis syn_module_defined=1 */ ;
    input \notGate[911]_keep ;
    output \notGate[912] ;
    
    wire \notGate[911]_keep  /* synthesis alspreserve=1 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(25[15:22])
    
    LUT4 I1 (.A(\notGate[911]_keep ), .B(\notGate[911]_keep ), .C(\notGate[911]_keep ), 
         .D(\notGate[911]_keep ), .Z(\notGate[912] )) /* synthesis syn_instantiated=1, lut_function=((!D !C !B !A)+(!D !C !B A)+(!D !C B !A)+(!D !C B A)+(!D C !B !A)+(!D C !B A)+(!D C B !A)+(!D C B A)), LSE_LINE_FILE_ID=3, LSE_LCOL=13, LSE_RCOL=44, LSE_LLINE=32, LSE_RLINE=32 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(11[2:53])
    defparam I1.init = 16'b0000000011111111;
    
endmodule
//
// Verilog Description of module inverter_U97
//

module inverter_U97 (\notGate[910]_keep , \notGate[911] ) /* synthesis syn_module_defined=1 */ ;
    input \notGate[910]_keep ;
    output \notGate[911] ;
    
    wire \notGate[910]_keep  /* synthesis alspreserve=1 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(25[15:22])
    
    LUT4 I1 (.A(\notGate[910]_keep ), .B(\notGate[910]_keep ), .C(\notGate[910]_keep ), 
         .D(\notGate[910]_keep ), .Z(\notGate[911] )) /* synthesis syn_instantiated=1, lut_function=((!D !C !B !A)+(!D !C !B A)+(!D !C B !A)+(!D !C B A)+(!D C !B !A)+(!D C !B A)+(!D C B !A)+(!D C B A)), LSE_LINE_FILE_ID=3, LSE_LCOL=13, LSE_RCOL=44, LSE_LLINE=32, LSE_RLINE=32 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(11[2:53])
    defparam I1.init = 16'b0000000011111111;
    
endmodule
//
// Verilog Description of module inverter_U98
//

module inverter_U98 (\notGate[909]_keep , \notGate[910] ) /* synthesis syn_module_defined=1 */ ;
    input \notGate[909]_keep ;
    output \notGate[910] ;
    
    wire \notGate[909]_keep  /* synthesis alspreserve=1 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(25[15:22])
    
    LUT4 I1 (.A(\notGate[909]_keep ), .B(\notGate[909]_keep ), .C(\notGate[909]_keep ), 
         .D(\notGate[909]_keep ), .Z(\notGate[910] )) /* synthesis syn_instantiated=1, lut_function=((!D !C !B !A)+(!D !C !B A)+(!D !C B !A)+(!D !C B A)+(!D C !B !A)+(!D C !B A)+(!D C B !A)+(!D C B A)), LSE_LINE_FILE_ID=3, LSE_LCOL=13, LSE_RCOL=44, LSE_LLINE=32, LSE_RLINE=32 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(11[2:53])
    defparam I1.init = 16'b0000000011111111;
    
endmodule
//
// Verilog Description of module inverter_U99
//

module inverter_U99 (\notGate[89]_keep , \notGate[90] ) /* synthesis syn_module_defined=1 */ ;
    input \notGate[89]_keep ;
    output \notGate[90] ;
    
    wire \notGate[89]_keep  /* synthesis alspreserve=1 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(25[15:22])
    
    LUT4 I1 (.A(\notGate[89]_keep ), .B(\notGate[89]_keep ), .C(\notGate[89]_keep ), 
         .D(\notGate[89]_keep ), .Z(\notGate[90] )) /* synthesis syn_instantiated=1, lut_function=((!D !C !B !A)+(!D !C !B A)+(!D !C B !A)+(!D !C B A)+(!D C !B !A)+(!D C !B A)+(!D C B !A)+(!D C B A)), LSE_LINE_FILE_ID=3, LSE_LCOL=13, LSE_RCOL=44, LSE_LLINE=32, LSE_RLINE=32 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(11[2:53])
    defparam I1.init = 16'b0000000011111111;
    
endmodule
//
// Verilog Description of module inverter_U100
//

module inverter_U100 (\notGate[908]_keep , \notGate[909] ) /* synthesis syn_module_defined=1 */ ;
    input \notGate[908]_keep ;
    output \notGate[909] ;
    
    wire \notGate[908]_keep  /* synthesis alspreserve=1 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(25[15:22])
    
    LUT4 I1 (.A(\notGate[908]_keep ), .B(\notGate[908]_keep ), .C(\notGate[908]_keep ), 
         .D(\notGate[908]_keep ), .Z(\notGate[909] )) /* synthesis syn_instantiated=1, lut_function=((!D !C !B !A)+(!D !C !B A)+(!D !C B !A)+(!D !C B A)+(!D C !B !A)+(!D C !B A)+(!D C B !A)+(!D C B A)), LSE_LINE_FILE_ID=3, LSE_LCOL=13, LSE_RCOL=44, LSE_LLINE=32, LSE_RLINE=32 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(11[2:53])
    defparam I1.init = 16'b0000000011111111;
    
endmodule
//
// Verilog Description of module inverter_U101
//

module inverter_U101 (\notGate[907]_keep , \notGate[908] ) /* synthesis syn_module_defined=1 */ ;
    input \notGate[907]_keep ;
    output \notGate[908] ;
    
    wire \notGate[907]_keep  /* synthesis alspreserve=1 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(25[15:22])
    
    LUT4 I1 (.A(\notGate[907]_keep ), .B(\notGate[907]_keep ), .C(\notGate[907]_keep ), 
         .D(\notGate[907]_keep ), .Z(\notGate[908] )) /* synthesis syn_instantiated=1, lut_function=((!D !C !B !A)+(!D !C !B A)+(!D !C B !A)+(!D !C B A)+(!D C !B !A)+(!D C !B A)+(!D C B !A)+(!D C B A)), LSE_LINE_FILE_ID=3, LSE_LCOL=13, LSE_RCOL=44, LSE_LLINE=32, LSE_RLINE=32 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(11[2:53])
    defparam I1.init = 16'b0000000011111111;
    
endmodule
//
// Verilog Description of module inverter_U102
//

module inverter_U102 (\notGate[906]_keep , \notGate[907] ) /* synthesis syn_module_defined=1 */ ;
    input \notGate[906]_keep ;
    output \notGate[907] ;
    
    wire \notGate[906]_keep  /* synthesis alspreserve=1 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(25[15:22])
    
    LUT4 I1 (.A(\notGate[906]_keep ), .B(\notGate[906]_keep ), .C(\notGate[906]_keep ), 
         .D(\notGate[906]_keep ), .Z(\notGate[907] )) /* synthesis syn_instantiated=1, lut_function=((!D !C !B !A)+(!D !C !B A)+(!D !C B !A)+(!D !C B A)+(!D C !B !A)+(!D C !B A)+(!D C B !A)+(!D C B A)), LSE_LINE_FILE_ID=3, LSE_LCOL=13, LSE_RCOL=44, LSE_LLINE=32, LSE_RLINE=32 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(11[2:53])
    defparam I1.init = 16'b0000000011111111;
    
endmodule
//
// Verilog Description of module inverter_U103
//

module inverter_U103 (\notGate[905]_keep , \notGate[906] ) /* synthesis syn_module_defined=1 */ ;
    input \notGate[905]_keep ;
    output \notGate[906] ;
    
    wire \notGate[905]_keep  /* synthesis alspreserve=1 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(25[15:22])
    
    LUT4 I1 (.A(\notGate[905]_keep ), .B(\notGate[905]_keep ), .C(\notGate[905]_keep ), 
         .D(\notGate[905]_keep ), .Z(\notGate[906] )) /* synthesis syn_instantiated=1, lut_function=((!D !C !B !A)+(!D !C !B A)+(!D !C B !A)+(!D !C B A)+(!D C !B !A)+(!D C !B A)+(!D C B !A)+(!D C B A)), LSE_LINE_FILE_ID=3, LSE_LCOL=13, LSE_RCOL=44, LSE_LLINE=32, LSE_RLINE=32 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(11[2:53])
    defparam I1.init = 16'b0000000011111111;
    
endmodule
//
// Verilog Description of module inverter_U104
//

module inverter_U104 (\notGate[904]_keep , \notGate[905] ) /* synthesis syn_module_defined=1 */ ;
    input \notGate[904]_keep ;
    output \notGate[905] ;
    
    wire \notGate[904]_keep  /* synthesis alspreserve=1 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(25[15:22])
    
    LUT4 I1 (.A(\notGate[904]_keep ), .B(\notGate[904]_keep ), .C(\notGate[904]_keep ), 
         .D(\notGate[904]_keep ), .Z(\notGate[905] )) /* synthesis syn_instantiated=1, lut_function=((!D !C !B !A)+(!D !C !B A)+(!D !C B !A)+(!D !C B A)+(!D C !B !A)+(!D C !B A)+(!D C B !A)+(!D C B A)), LSE_LINE_FILE_ID=3, LSE_LCOL=13, LSE_RCOL=44, LSE_LLINE=32, LSE_RLINE=32 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(11[2:53])
    defparam I1.init = 16'b0000000011111111;
    
endmodule
//
// Verilog Description of module inverter_U105
//

module inverter_U105 (\notGate[903]_keep , \notGate[904] ) /* synthesis syn_module_defined=1 */ ;
    input \notGate[903]_keep ;
    output \notGate[904] ;
    
    wire \notGate[903]_keep  /* synthesis alspreserve=1 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(25[15:22])
    
    LUT4 I1 (.A(\notGate[903]_keep ), .B(\notGate[903]_keep ), .C(\notGate[903]_keep ), 
         .D(\notGate[903]_keep ), .Z(\notGate[904] )) /* synthesis syn_instantiated=1, lut_function=((!D !C !B !A)+(!D !C !B A)+(!D !C B !A)+(!D !C B A)+(!D C !B !A)+(!D C !B A)+(!D C B !A)+(!D C B A)), LSE_LINE_FILE_ID=3, LSE_LCOL=13, LSE_RCOL=44, LSE_LLINE=32, LSE_RLINE=32 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(11[2:53])
    defparam I1.init = 16'b0000000011111111;
    
endmodule
//
// Verilog Description of module inverter_U106
//

module inverter_U106 (\notGate[902]_keep , \notGate[903] ) /* synthesis syn_module_defined=1 */ ;
    input \notGate[902]_keep ;
    output \notGate[903] ;
    
    wire \notGate[902]_keep  /* synthesis alspreserve=1 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(25[15:22])
    
    LUT4 I1 (.A(\notGate[902]_keep ), .B(\notGate[902]_keep ), .C(\notGate[902]_keep ), 
         .D(\notGate[902]_keep ), .Z(\notGate[903] )) /* synthesis syn_instantiated=1, lut_function=((!D !C !B !A)+(!D !C !B A)+(!D !C B !A)+(!D !C B A)+(!D C !B !A)+(!D C !B A)+(!D C B !A)+(!D C B A)), LSE_LINE_FILE_ID=3, LSE_LCOL=13, LSE_RCOL=44, LSE_LLINE=32, LSE_RLINE=32 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(11[2:53])
    defparam I1.init = 16'b0000000011111111;
    
endmodule
//
// Verilog Description of module inverter_U107
//

module inverter_U107 (\notGate[901]_keep , \notGate[902] ) /* synthesis syn_module_defined=1 */ ;
    input \notGate[901]_keep ;
    output \notGate[902] ;
    
    wire \notGate[901]_keep  /* synthesis alspreserve=1 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(25[15:22])
    
    LUT4 I1 (.A(\notGate[901]_keep ), .B(\notGate[901]_keep ), .C(\notGate[901]_keep ), 
         .D(\notGate[901]_keep ), .Z(\notGate[902] )) /* synthesis syn_instantiated=1, lut_function=((!D !C !B !A)+(!D !C !B A)+(!D !C B !A)+(!D !C B A)+(!D C !B !A)+(!D C !B A)+(!D C B !A)+(!D C B A)), LSE_LINE_FILE_ID=3, LSE_LCOL=13, LSE_RCOL=44, LSE_LLINE=32, LSE_RLINE=32 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(11[2:53])
    defparam I1.init = 16'b0000000011111111;
    
endmodule
//
// Verilog Description of module inverter_U108
//

module inverter_U108 (\notGate[900]_keep , \notGate[901] ) /* synthesis syn_module_defined=1 */ ;
    input \notGate[900]_keep ;
    output \notGate[901] ;
    
    wire \notGate[900]_keep  /* synthesis alspreserve=1 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(25[15:22])
    
    LUT4 I1 (.A(\notGate[900]_keep ), .B(\notGate[900]_keep ), .C(\notGate[900]_keep ), 
         .D(\notGate[900]_keep ), .Z(\notGate[901] )) /* synthesis syn_instantiated=1, lut_function=((!D !C !B !A)+(!D !C !B A)+(!D !C B !A)+(!D !C B A)+(!D C !B !A)+(!D C !B A)+(!D C B !A)+(!D C B A)), LSE_LINE_FILE_ID=3, LSE_LCOL=13, LSE_RCOL=44, LSE_LLINE=32, LSE_RLINE=32 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(11[2:53])
    defparam I1.init = 16'b0000000011111111;
    
endmodule
//
// Verilog Description of module inverter_U109
//

module inverter_U109 (\notGate[899]_keep , \notGate[900] ) /* synthesis syn_module_defined=1 */ ;
    input \notGate[899]_keep ;
    output \notGate[900] ;
    
    wire \notGate[899]_keep  /* synthesis alspreserve=1 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(25[15:22])
    
    LUT4 I1 (.A(\notGate[899]_keep ), .B(\notGate[899]_keep ), .C(\notGate[899]_keep ), 
         .D(\notGate[899]_keep ), .Z(\notGate[900] )) /* synthesis syn_instantiated=1, lut_function=((!D !C !B !A)+(!D !C !B A)+(!D !C B !A)+(!D !C B A)+(!D C !B !A)+(!D C !B A)+(!D C B !A)+(!D C B A)), LSE_LINE_FILE_ID=3, LSE_LCOL=13, LSE_RCOL=44, LSE_LLINE=32, LSE_RLINE=32 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(11[2:53])
    defparam I1.init = 16'b0000000011111111;
    
endmodule
//
// Verilog Description of module inverter_U110
//

module inverter_U110 (\notGate[7]_keep , \notGate[8] ) /* synthesis syn_module_defined=1 */ ;
    input \notGate[7]_keep ;
    output \notGate[8] ;
    
    wire \notGate[7]_keep  /* synthesis alspreserve=1 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(25[15:22])
    
    LUT4 I1 (.A(\notGate[7]_keep ), .B(\notGate[7]_keep ), .C(\notGate[7]_keep ), 
         .D(\notGate[7]_keep ), .Z(\notGate[8] )) /* synthesis syn_instantiated=1, lut_function=((!D !C !B !A)+(!D !C !B A)+(!D !C B !A)+(!D !C B A)+(!D C !B !A)+(!D C !B A)+(!D C B !A)+(!D C B A)), LSE_LINE_FILE_ID=3, LSE_LCOL=13, LSE_RCOL=44, LSE_LLINE=32, LSE_RLINE=32 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(11[2:53])
    defparam I1.init = 16'b0000000011111111;
    
endmodule
//
// Verilog Description of module inverter_U111
//

module inverter_U111 (\notGate[88]_keep , \notGate[89] ) /* synthesis syn_module_defined=1 */ ;
    input \notGate[88]_keep ;
    output \notGate[89] ;
    
    wire \notGate[88]_keep  /* synthesis alspreserve=1 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(25[15:22])
    
    LUT4 I1 (.A(\notGate[88]_keep ), .B(\notGate[88]_keep ), .C(\notGate[88]_keep ), 
         .D(\notGate[88]_keep ), .Z(\notGate[89] )) /* synthesis syn_instantiated=1, lut_function=((!D !C !B !A)+(!D !C !B A)+(!D !C B !A)+(!D !C B A)+(!D C !B !A)+(!D C !B A)+(!D C B !A)+(!D C B A)), LSE_LINE_FILE_ID=3, LSE_LCOL=13, LSE_RCOL=44, LSE_LLINE=32, LSE_RLINE=32 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(11[2:53])
    defparam I1.init = 16'b0000000011111111;
    
endmodule
//
// Verilog Description of module inverter_U112
//

module inverter_U112 (\notGate[898]_keep , \notGate[899] ) /* synthesis syn_module_defined=1 */ ;
    input \notGate[898]_keep ;
    output \notGate[899] ;
    
    wire \notGate[898]_keep  /* synthesis alspreserve=1 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(25[15:22])
    
    LUT4 I1 (.A(\notGate[898]_keep ), .B(\notGate[898]_keep ), .C(\notGate[898]_keep ), 
         .D(\notGate[898]_keep ), .Z(\notGate[899] )) /* synthesis syn_instantiated=1, lut_function=((!D !C !B !A)+(!D !C !B A)+(!D !C B !A)+(!D !C B A)+(!D C !B !A)+(!D C !B A)+(!D C B !A)+(!D C B A)), LSE_LINE_FILE_ID=3, LSE_LCOL=13, LSE_RCOL=44, LSE_LLINE=32, LSE_RLINE=32 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(11[2:53])
    defparam I1.init = 16'b0000000011111111;
    
endmodule
//
// Verilog Description of module inverter_U113
//

module inverter_U113 (\notGate[897]_keep , \notGate[898] ) /* synthesis syn_module_defined=1 */ ;
    input \notGate[897]_keep ;
    output \notGate[898] ;
    
    wire \notGate[897]_keep  /* synthesis alspreserve=1 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(25[15:22])
    
    LUT4 I1 (.A(\notGate[897]_keep ), .B(\notGate[897]_keep ), .C(\notGate[897]_keep ), 
         .D(\notGate[897]_keep ), .Z(\notGate[898] )) /* synthesis syn_instantiated=1, lut_function=((!D !C !B !A)+(!D !C !B A)+(!D !C B !A)+(!D !C B A)+(!D C !B !A)+(!D C !B A)+(!D C B !A)+(!D C B A)), LSE_LINE_FILE_ID=3, LSE_LCOL=13, LSE_RCOL=44, LSE_LLINE=32, LSE_RLINE=32 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(11[2:53])
    defparam I1.init = 16'b0000000011111111;
    
endmodule
//
// Verilog Description of module inverter_U114
//

module inverter_U114 (\notGate[896]_keep , \notGate[897] ) /* synthesis syn_module_defined=1 */ ;
    input \notGate[896]_keep ;
    output \notGate[897] ;
    
    wire \notGate[896]_keep  /* synthesis alspreserve=1 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(25[15:22])
    
    LUT4 I1 (.A(\notGate[896]_keep ), .B(\notGate[896]_keep ), .C(\notGate[896]_keep ), 
         .D(\notGate[896]_keep ), .Z(\notGate[897] )) /* synthesis syn_instantiated=1, lut_function=((!D !C !B !A)+(!D !C !B A)+(!D !C B !A)+(!D !C B A)+(!D C !B !A)+(!D C !B A)+(!D C B !A)+(!D C B A)), LSE_LINE_FILE_ID=3, LSE_LCOL=13, LSE_RCOL=44, LSE_LLINE=32, LSE_RLINE=32 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(11[2:53])
    defparam I1.init = 16'b0000000011111111;
    
endmodule
//
// Verilog Description of module inverter_U115
//

module inverter_U115 (\notGate[895]_keep , \notGate[896] ) /* synthesis syn_module_defined=1 */ ;
    input \notGate[895]_keep ;
    output \notGate[896] ;
    
    wire \notGate[895]_keep  /* synthesis alspreserve=1 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(25[15:22])
    
    LUT4 I1 (.A(\notGate[895]_keep ), .B(\notGate[895]_keep ), .C(\notGate[895]_keep ), 
         .D(\notGate[895]_keep ), .Z(\notGate[896] )) /* synthesis syn_instantiated=1, lut_function=((!D !C !B !A)+(!D !C !B A)+(!D !C B !A)+(!D !C B A)+(!D C !B !A)+(!D C !B A)+(!D C B !A)+(!D C B A)), LSE_LINE_FILE_ID=3, LSE_LCOL=13, LSE_RCOL=44, LSE_LLINE=32, LSE_RLINE=32 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(11[2:53])
    defparam I1.init = 16'b0000000011111111;
    
endmodule
//
// Verilog Description of module inverter_U116
//

module inverter_U116 (\notGate[894]_keep , \notGate[895] ) /* synthesis syn_module_defined=1 */ ;
    input \notGate[894]_keep ;
    output \notGate[895] ;
    
    wire \notGate[894]_keep  /* synthesis alspreserve=1 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(25[15:22])
    
    LUT4 I1 (.A(\notGate[894]_keep ), .B(\notGate[894]_keep ), .C(\notGate[894]_keep ), 
         .D(\notGate[894]_keep ), .Z(\notGate[895] )) /* synthesis syn_instantiated=1, lut_function=((!D !C !B !A)+(!D !C !B A)+(!D !C B !A)+(!D !C B A)+(!D C !B !A)+(!D C !B A)+(!D C B !A)+(!D C B A)), LSE_LINE_FILE_ID=3, LSE_LCOL=13, LSE_RCOL=44, LSE_LLINE=32, LSE_RLINE=32 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(11[2:53])
    defparam I1.init = 16'b0000000011111111;
    
endmodule
//
// Verilog Description of module inverter_U117
//

module inverter_U117 (\notGate[893]_keep , \notGate[894] ) /* synthesis syn_module_defined=1 */ ;
    input \notGate[893]_keep ;
    output \notGate[894] ;
    
    wire \notGate[893]_keep  /* synthesis alspreserve=1 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(25[15:22])
    
    LUT4 I1 (.A(\notGate[893]_keep ), .B(\notGate[893]_keep ), .C(\notGate[893]_keep ), 
         .D(\notGate[893]_keep ), .Z(\notGate[894] )) /* synthesis syn_instantiated=1, lut_function=((!D !C !B !A)+(!D !C !B A)+(!D !C B !A)+(!D !C B A)+(!D C !B !A)+(!D C !B A)+(!D C B !A)+(!D C B A)), LSE_LINE_FILE_ID=3, LSE_LCOL=13, LSE_RCOL=44, LSE_LLINE=32, LSE_RLINE=32 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(11[2:53])
    defparam I1.init = 16'b0000000011111111;
    
endmodule
//
// Verilog Description of module inverter_U118
//

module inverter_U118 (\notGate[892]_keep , \notGate[893] ) /* synthesis syn_module_defined=1 */ ;
    input \notGate[892]_keep ;
    output \notGate[893] ;
    
    wire \notGate[892]_keep  /* synthesis alspreserve=1 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(25[15:22])
    
    LUT4 I1 (.A(\notGate[892]_keep ), .B(\notGate[892]_keep ), .C(\notGate[892]_keep ), 
         .D(\notGate[892]_keep ), .Z(\notGate[893] )) /* synthesis syn_instantiated=1, lut_function=((!D !C !B !A)+(!D !C !B A)+(!D !C B !A)+(!D !C B A)+(!D C !B !A)+(!D C !B A)+(!D C B !A)+(!D C B A)), LSE_LINE_FILE_ID=3, LSE_LCOL=13, LSE_RCOL=44, LSE_LLINE=32, LSE_RLINE=32 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(11[2:53])
    defparam I1.init = 16'b0000000011111111;
    
endmodule
//
// Verilog Description of module inverter_U119
//

module inverter_U119 (\notGate[891]_keep , \notGate[892] ) /* synthesis syn_module_defined=1 */ ;
    input \notGate[891]_keep ;
    output \notGate[892] ;
    
    wire \notGate[891]_keep  /* synthesis alspreserve=1 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(25[15:22])
    
    LUT4 I1 (.A(\notGate[891]_keep ), .B(\notGate[891]_keep ), .C(\notGate[891]_keep ), 
         .D(\notGate[891]_keep ), .Z(\notGate[892] )) /* synthesis syn_instantiated=1, lut_function=((!D !C !B !A)+(!D !C !B A)+(!D !C B !A)+(!D !C B A)+(!D C !B !A)+(!D C !B A)+(!D C B !A)+(!D C B A)), LSE_LINE_FILE_ID=3, LSE_LCOL=13, LSE_RCOL=44, LSE_LLINE=32, LSE_RLINE=32 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(11[2:53])
    defparam I1.init = 16'b0000000011111111;
    
endmodule
//
// Verilog Description of module inverter_U120
//

module inverter_U120 (\notGate[890]_keep , \notGate[891] ) /* synthesis syn_module_defined=1 */ ;
    input \notGate[890]_keep ;
    output \notGate[891] ;
    
    wire \notGate[890]_keep  /* synthesis alspreserve=1 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(25[15:22])
    
    LUT4 I1 (.A(\notGate[890]_keep ), .B(\notGate[890]_keep ), .C(\notGate[890]_keep ), 
         .D(\notGate[890]_keep ), .Z(\notGate[891] )) /* synthesis syn_instantiated=1, lut_function=((!D !C !B !A)+(!D !C !B A)+(!D !C B !A)+(!D !C B A)+(!D C !B !A)+(!D C !B A)+(!D C B !A)+(!D C B A)), LSE_LINE_FILE_ID=3, LSE_LCOL=13, LSE_RCOL=44, LSE_LLINE=32, LSE_RLINE=32 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(11[2:53])
    defparam I1.init = 16'b0000000011111111;
    
endmodule
//
// Verilog Description of module inverter_U121
//

module inverter_U121 (\notGate[889]_keep , \notGate[890] ) /* synthesis syn_module_defined=1 */ ;
    input \notGate[889]_keep ;
    output \notGate[890] ;
    
    wire \notGate[889]_keep  /* synthesis alspreserve=1 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(25[15:22])
    
    LUT4 I1 (.A(\notGate[889]_keep ), .B(\notGate[889]_keep ), .C(\notGate[889]_keep ), 
         .D(\notGate[889]_keep ), .Z(\notGate[890] )) /* synthesis syn_instantiated=1, lut_function=((!D !C !B !A)+(!D !C !B A)+(!D !C B !A)+(!D !C B A)+(!D C !B !A)+(!D C !B A)+(!D C B !A)+(!D C B A)), LSE_LINE_FILE_ID=3, LSE_LCOL=13, LSE_RCOL=44, LSE_LLINE=32, LSE_RLINE=32 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(11[2:53])
    defparam I1.init = 16'b0000000011111111;
    
endmodule
//
// Verilog Description of module inverter_U122
//

module inverter_U122 (\notGate[87]_keep , \notGate[88] ) /* synthesis syn_module_defined=1 */ ;
    input \notGate[87]_keep ;
    output \notGate[88] ;
    
    wire \notGate[87]_keep  /* synthesis alspreserve=1 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(25[15:22])
    
    LUT4 I1 (.A(\notGate[87]_keep ), .B(\notGate[87]_keep ), .C(\notGate[87]_keep ), 
         .D(\notGate[87]_keep ), .Z(\notGate[88] )) /* synthesis syn_instantiated=1, lut_function=((!D !C !B !A)+(!D !C !B A)+(!D !C B !A)+(!D !C B A)+(!D C !B !A)+(!D C !B A)+(!D C B !A)+(!D C B A)), LSE_LINE_FILE_ID=3, LSE_LCOL=13, LSE_RCOL=44, LSE_LLINE=32, LSE_RLINE=32 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(11[2:53])
    defparam I1.init = 16'b0000000011111111;
    
endmodule
//
// Verilog Description of module inverter_U123
//

module inverter_U123 (\notGate[888]_keep , \notGate[889] ) /* synthesis syn_module_defined=1 */ ;
    input \notGate[888]_keep ;
    output \notGate[889] ;
    
    wire \notGate[888]_keep  /* synthesis alspreserve=1 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(25[15:22])
    
    LUT4 I1 (.A(\notGate[888]_keep ), .B(\notGate[888]_keep ), .C(\notGate[888]_keep ), 
         .D(\notGate[888]_keep ), .Z(\notGate[889] )) /* synthesis syn_instantiated=1, lut_function=((!D !C !B !A)+(!D !C !B A)+(!D !C B !A)+(!D !C B A)+(!D C !B !A)+(!D C !B A)+(!D C B !A)+(!D C B A)), LSE_LINE_FILE_ID=3, LSE_LCOL=13, LSE_RCOL=44, LSE_LLINE=32, LSE_RLINE=32 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(11[2:53])
    defparam I1.init = 16'b0000000011111111;
    
endmodule
//
// Verilog Description of module inverter_U124
//

module inverter_U124 (\notGate[887]_keep , \notGate[888] ) /* synthesis syn_module_defined=1 */ ;
    input \notGate[887]_keep ;
    output \notGate[888] ;
    
    wire \notGate[887]_keep  /* synthesis alspreserve=1 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(25[15:22])
    
    LUT4 I1 (.A(\notGate[887]_keep ), .B(\notGate[887]_keep ), .C(\notGate[887]_keep ), 
         .D(\notGate[887]_keep ), .Z(\notGate[888] )) /* synthesis syn_instantiated=1, lut_function=((!D !C !B !A)+(!D !C !B A)+(!D !C B !A)+(!D !C B A)+(!D C !B !A)+(!D C !B A)+(!D C B !A)+(!D C B A)), LSE_LINE_FILE_ID=3, LSE_LCOL=13, LSE_RCOL=44, LSE_LLINE=32, LSE_RLINE=32 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(11[2:53])
    defparam I1.init = 16'b0000000011111111;
    
endmodule
//
// Verilog Description of module inverter_U125
//

module inverter_U125 (\notGate[886]_keep , \notGate[887] ) /* synthesis syn_module_defined=1 */ ;
    input \notGate[886]_keep ;
    output \notGate[887] ;
    
    wire \notGate[886]_keep  /* synthesis alspreserve=1 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(25[15:22])
    
    LUT4 I1 (.A(\notGate[886]_keep ), .B(\notGate[886]_keep ), .C(\notGate[886]_keep ), 
         .D(\notGate[886]_keep ), .Z(\notGate[887] )) /* synthesis syn_instantiated=1, lut_function=((!D !C !B !A)+(!D !C !B A)+(!D !C B !A)+(!D !C B A)+(!D C !B !A)+(!D C !B A)+(!D C B !A)+(!D C B A)), LSE_LINE_FILE_ID=3, LSE_LCOL=13, LSE_RCOL=44, LSE_LLINE=32, LSE_RLINE=32 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(11[2:53])
    defparam I1.init = 16'b0000000011111111;
    
endmodule
//
// Verilog Description of module inverter_U126
//

module inverter_U126 (\notGate[885]_keep , \notGate[886] ) /* synthesis syn_module_defined=1 */ ;
    input \notGate[885]_keep ;
    output \notGate[886] ;
    
    wire \notGate[885]_keep  /* synthesis alspreserve=1 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(25[15:22])
    
    LUT4 I1 (.A(\notGate[885]_keep ), .B(\notGate[885]_keep ), .C(\notGate[885]_keep ), 
         .D(\notGate[885]_keep ), .Z(\notGate[886] )) /* synthesis syn_instantiated=1, lut_function=((!D !C !B !A)+(!D !C !B A)+(!D !C B !A)+(!D !C B A)+(!D C !B !A)+(!D C !B A)+(!D C B !A)+(!D C B A)), LSE_LINE_FILE_ID=3, LSE_LCOL=13, LSE_RCOL=44, LSE_LLINE=32, LSE_RLINE=32 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(11[2:53])
    defparam I1.init = 16'b0000000011111111;
    
endmodule
//
// Verilog Description of module inverter_U127
//

module inverter_U127 (\notGate[884]_keep , \notGate[885] ) /* synthesis syn_module_defined=1 */ ;
    input \notGate[884]_keep ;
    output \notGate[885] ;
    
    wire \notGate[884]_keep  /* synthesis alspreserve=1 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(25[15:22])
    
    LUT4 I1 (.A(\notGate[884]_keep ), .B(\notGate[884]_keep ), .C(\notGate[884]_keep ), 
         .D(\notGate[884]_keep ), .Z(\notGate[885] )) /* synthesis syn_instantiated=1, lut_function=((!D !C !B !A)+(!D !C !B A)+(!D !C B !A)+(!D !C B A)+(!D C !B !A)+(!D C !B A)+(!D C B !A)+(!D C B A)), LSE_LINE_FILE_ID=3, LSE_LCOL=13, LSE_RCOL=44, LSE_LLINE=32, LSE_RLINE=32 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(11[2:53])
    defparam I1.init = 16'b0000000011111111;
    
endmodule
//
// Verilog Description of module inverter_U128
//

module inverter_U128 (\notGate[883]_keep , \notGate[884] ) /* synthesis syn_module_defined=1 */ ;
    input \notGate[883]_keep ;
    output \notGate[884] ;
    
    wire \notGate[883]_keep  /* synthesis alspreserve=1 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(25[15:22])
    
    LUT4 I1 (.A(\notGate[883]_keep ), .B(\notGate[883]_keep ), .C(\notGate[883]_keep ), 
         .D(\notGate[883]_keep ), .Z(\notGate[884] )) /* synthesis syn_instantiated=1, lut_function=((!D !C !B !A)+(!D !C !B A)+(!D !C B !A)+(!D !C B A)+(!D C !B !A)+(!D C !B A)+(!D C B !A)+(!D C B A)), LSE_LINE_FILE_ID=3, LSE_LCOL=13, LSE_RCOL=44, LSE_LLINE=32, LSE_RLINE=32 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(11[2:53])
    defparam I1.init = 16'b0000000011111111;
    
endmodule
//
// Verilog Description of module inverter_U129
//

module inverter_U129 (\notGate[882]_keep , \notGate[883] ) /* synthesis syn_module_defined=1 */ ;
    input \notGate[882]_keep ;
    output \notGate[883] ;
    
    wire \notGate[882]_keep  /* synthesis alspreserve=1 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(25[15:22])
    
    LUT4 I1 (.A(\notGate[882]_keep ), .B(\notGate[882]_keep ), .C(\notGate[882]_keep ), 
         .D(\notGate[882]_keep ), .Z(\notGate[883] )) /* synthesis syn_instantiated=1, lut_function=((!D !C !B !A)+(!D !C !B A)+(!D !C B !A)+(!D !C B A)+(!D C !B !A)+(!D C !B A)+(!D C B !A)+(!D C B A)), LSE_LINE_FILE_ID=3, LSE_LCOL=13, LSE_RCOL=44, LSE_LLINE=32, LSE_RLINE=32 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(11[2:53])
    defparam I1.init = 16'b0000000011111111;
    
endmodule
//
// Verilog Description of module inverter_U130
//

module inverter_U130 (\notGate[881]_keep , \notGate[882] ) /* synthesis syn_module_defined=1 */ ;
    input \notGate[881]_keep ;
    output \notGate[882] ;
    
    wire \notGate[881]_keep  /* synthesis alspreserve=1 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(25[15:22])
    
    LUT4 I1 (.A(\notGate[881]_keep ), .B(\notGate[881]_keep ), .C(\notGate[881]_keep ), 
         .D(\notGate[881]_keep ), .Z(\notGate[882] )) /* synthesis syn_instantiated=1, lut_function=((!D !C !B !A)+(!D !C !B A)+(!D !C B !A)+(!D !C B A)+(!D C !B !A)+(!D C !B A)+(!D C B !A)+(!D C B A)), LSE_LINE_FILE_ID=3, LSE_LCOL=13, LSE_RCOL=44, LSE_LLINE=32, LSE_RLINE=32 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(11[2:53])
    defparam I1.init = 16'b0000000011111111;
    
endmodule
//
// Verilog Description of module inverter_U131
//

module inverter_U131 (\notGate[880]_keep , \notGate[881] ) /* synthesis syn_module_defined=1 */ ;
    input \notGate[880]_keep ;
    output \notGate[881] ;
    
    wire \notGate[880]_keep  /* synthesis alspreserve=1 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(25[15:22])
    
    LUT4 I1 (.A(\notGate[880]_keep ), .B(\notGate[880]_keep ), .C(\notGate[880]_keep ), 
         .D(\notGate[880]_keep ), .Z(\notGate[881] )) /* synthesis syn_instantiated=1, lut_function=((!D !C !B !A)+(!D !C !B A)+(!D !C B !A)+(!D !C B A)+(!D C !B !A)+(!D C !B A)+(!D C B !A)+(!D C B A)), LSE_LINE_FILE_ID=3, LSE_LCOL=13, LSE_RCOL=44, LSE_LLINE=32, LSE_RLINE=32 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(11[2:53])
    defparam I1.init = 16'b0000000011111111;
    
endmodule
//
// Verilog Description of module inverter_U132
//

module inverter_U132 (\notGate[879]_keep , \notGate[880] ) /* synthesis syn_module_defined=1 */ ;
    input \notGate[879]_keep ;
    output \notGate[880] ;
    
    wire \notGate[879]_keep  /* synthesis alspreserve=1 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(25[15:22])
    
    LUT4 I1 (.A(\notGate[879]_keep ), .B(\notGate[879]_keep ), .C(\notGate[879]_keep ), 
         .D(\notGate[879]_keep ), .Z(\notGate[880] )) /* synthesis syn_instantiated=1, lut_function=((!D !C !B !A)+(!D !C !B A)+(!D !C B !A)+(!D !C B A)+(!D C !B !A)+(!D C !B A)+(!D C B !A)+(!D C B A)), LSE_LINE_FILE_ID=3, LSE_LCOL=13, LSE_RCOL=44, LSE_LLINE=32, LSE_RLINE=32 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(11[2:53])
    defparam I1.init = 16'b0000000011111111;
    
endmodule
//
// Verilog Description of module inverter_U133
//

module inverter_U133 (\notGate[86]_keep , \notGate[87] ) /* synthesis syn_module_defined=1 */ ;
    input \notGate[86]_keep ;
    output \notGate[87] ;
    
    wire \notGate[86]_keep  /* synthesis alspreserve=1 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(25[15:22])
    
    LUT4 I1 (.A(\notGate[86]_keep ), .B(\notGate[86]_keep ), .C(\notGate[86]_keep ), 
         .D(\notGate[86]_keep ), .Z(\notGate[87] )) /* synthesis syn_instantiated=1, lut_function=((!D !C !B !A)+(!D !C !B A)+(!D !C B !A)+(!D !C B A)+(!D C !B !A)+(!D C !B A)+(!D C B !A)+(!D C B A)), LSE_LINE_FILE_ID=3, LSE_LCOL=13, LSE_RCOL=44, LSE_LLINE=32, LSE_RLINE=32 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(11[2:53])
    defparam I1.init = 16'b0000000011111111;
    
endmodule
//
// Verilog Description of module inverter_U134
//

module inverter_U134 (\notGate[878]_keep , \notGate[879] ) /* synthesis syn_module_defined=1 */ ;
    input \notGate[878]_keep ;
    output \notGate[879] ;
    
    wire \notGate[878]_keep  /* synthesis alspreserve=1 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(25[15:22])
    
    LUT4 I1 (.A(\notGate[878]_keep ), .B(\notGate[878]_keep ), .C(\notGate[878]_keep ), 
         .D(\notGate[878]_keep ), .Z(\notGate[879] )) /* synthesis syn_instantiated=1, lut_function=((!D !C !B !A)+(!D !C !B A)+(!D !C B !A)+(!D !C B A)+(!D C !B !A)+(!D C !B A)+(!D C B !A)+(!D C B A)), LSE_LINE_FILE_ID=3, LSE_LCOL=13, LSE_RCOL=44, LSE_LLINE=32, LSE_RLINE=32 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(11[2:53])
    defparam I1.init = 16'b0000000011111111;
    
endmodule
//
// Verilog Description of module inverter_U135
//

module inverter_U135 (\notGate[877]_keep , \notGate[878] ) /* synthesis syn_module_defined=1 */ ;
    input \notGate[877]_keep ;
    output \notGate[878] ;
    
    wire \notGate[877]_keep  /* synthesis alspreserve=1 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(25[15:22])
    
    LUT4 I1 (.A(\notGate[877]_keep ), .B(\notGate[877]_keep ), .C(\notGate[877]_keep ), 
         .D(\notGate[877]_keep ), .Z(\notGate[878] )) /* synthesis syn_instantiated=1, lut_function=((!D !C !B !A)+(!D !C !B A)+(!D !C B !A)+(!D !C B A)+(!D C !B !A)+(!D C !B A)+(!D C B !A)+(!D C B A)), LSE_LINE_FILE_ID=3, LSE_LCOL=13, LSE_RCOL=44, LSE_LLINE=32, LSE_RLINE=32 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(11[2:53])
    defparam I1.init = 16'b0000000011111111;
    
endmodule
//
// Verilog Description of module inverter_U136
//

module inverter_U136 (\notGate[876]_keep , \notGate[877] ) /* synthesis syn_module_defined=1 */ ;
    input \notGate[876]_keep ;
    output \notGate[877] ;
    
    wire \notGate[876]_keep  /* synthesis alspreserve=1 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(25[15:22])
    
    LUT4 I1 (.A(\notGate[876]_keep ), .B(\notGate[876]_keep ), .C(\notGate[876]_keep ), 
         .D(\notGate[876]_keep ), .Z(\notGate[877] )) /* synthesis syn_instantiated=1, lut_function=((!D !C !B !A)+(!D !C !B A)+(!D !C B !A)+(!D !C B A)+(!D C !B !A)+(!D C !B A)+(!D C B !A)+(!D C B A)), LSE_LINE_FILE_ID=3, LSE_LCOL=13, LSE_RCOL=44, LSE_LLINE=32, LSE_RLINE=32 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(11[2:53])
    defparam I1.init = 16'b0000000011111111;
    
endmodule
//
// Verilog Description of module inverter_U137
//

module inverter_U137 (\notGate[875]_keep , \notGate[876] ) /* synthesis syn_module_defined=1 */ ;
    input \notGate[875]_keep ;
    output \notGate[876] ;
    
    wire \notGate[875]_keep  /* synthesis alspreserve=1 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(25[15:22])
    
    LUT4 I1 (.A(\notGate[875]_keep ), .B(\notGate[875]_keep ), .C(\notGate[875]_keep ), 
         .D(\notGate[875]_keep ), .Z(\notGate[876] )) /* synthesis syn_instantiated=1, lut_function=((!D !C !B !A)+(!D !C !B A)+(!D !C B !A)+(!D !C B A)+(!D C !B !A)+(!D C !B A)+(!D C B !A)+(!D C B A)), LSE_LINE_FILE_ID=3, LSE_LCOL=13, LSE_RCOL=44, LSE_LLINE=32, LSE_RLINE=32 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(11[2:53])
    defparam I1.init = 16'b0000000011111111;
    
endmodule
//
// Verilog Description of module inverter_U138
//

module inverter_U138 (\notGate[874]_keep , \notGate[875] ) /* synthesis syn_module_defined=1 */ ;
    input \notGate[874]_keep ;
    output \notGate[875] ;
    
    wire \notGate[874]_keep  /* synthesis alspreserve=1 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(25[15:22])
    
    LUT4 I1 (.A(\notGate[874]_keep ), .B(\notGate[874]_keep ), .C(\notGate[874]_keep ), 
         .D(\notGate[874]_keep ), .Z(\notGate[875] )) /* synthesis syn_instantiated=1, lut_function=((!D !C !B !A)+(!D !C !B A)+(!D !C B !A)+(!D !C B A)+(!D C !B !A)+(!D C !B A)+(!D C B !A)+(!D C B A)), LSE_LINE_FILE_ID=3, LSE_LCOL=13, LSE_RCOL=44, LSE_LLINE=32, LSE_RLINE=32 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(11[2:53])
    defparam I1.init = 16'b0000000011111111;
    
endmodule
//
// Verilog Description of module inverter_U139
//

module inverter_U139 (\notGate[873]_keep , \notGate[874] ) /* synthesis syn_module_defined=1 */ ;
    input \notGate[873]_keep ;
    output \notGate[874] ;
    
    wire \notGate[873]_keep  /* synthesis alspreserve=1 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(25[15:22])
    
    LUT4 I1 (.A(\notGate[873]_keep ), .B(\notGate[873]_keep ), .C(\notGate[873]_keep ), 
         .D(\notGate[873]_keep ), .Z(\notGate[874] )) /* synthesis syn_instantiated=1, lut_function=((!D !C !B !A)+(!D !C !B A)+(!D !C B !A)+(!D !C B A)+(!D C !B !A)+(!D C !B A)+(!D C B !A)+(!D C B A)), LSE_LINE_FILE_ID=3, LSE_LCOL=13, LSE_RCOL=44, LSE_LLINE=32, LSE_RLINE=32 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(11[2:53])
    defparam I1.init = 16'b0000000011111111;
    
endmodule
//
// Verilog Description of module inverter_U140
//

module inverter_U140 (\notGate[872]_keep , \notGate[873] ) /* synthesis syn_module_defined=1 */ ;
    input \notGate[872]_keep ;
    output \notGate[873] ;
    
    wire \notGate[872]_keep  /* synthesis alspreserve=1 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(25[15:22])
    
    LUT4 I1 (.A(\notGate[872]_keep ), .B(\notGate[872]_keep ), .C(\notGate[872]_keep ), 
         .D(\notGate[872]_keep ), .Z(\notGate[873] )) /* synthesis syn_instantiated=1, lut_function=((!D !C !B !A)+(!D !C !B A)+(!D !C B !A)+(!D !C B A)+(!D C !B !A)+(!D C !B A)+(!D C B !A)+(!D C B A)), LSE_LINE_FILE_ID=3, LSE_LCOL=13, LSE_RCOL=44, LSE_LLINE=32, LSE_RLINE=32 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(11[2:53])
    defparam I1.init = 16'b0000000011111111;
    
endmodule
//
// Verilog Description of module inverter_U141
//

module inverter_U141 (\notGate[871]_keep , \notGate[872] ) /* synthesis syn_module_defined=1 */ ;
    input \notGate[871]_keep ;
    output \notGate[872] ;
    
    wire \notGate[871]_keep  /* synthesis alspreserve=1 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(25[15:22])
    
    LUT4 I1 (.A(\notGate[871]_keep ), .B(\notGate[871]_keep ), .C(\notGate[871]_keep ), 
         .D(\notGate[871]_keep ), .Z(\notGate[872] )) /* synthesis syn_instantiated=1, lut_function=((!D !C !B !A)+(!D !C !B A)+(!D !C B !A)+(!D !C B A)+(!D C !B !A)+(!D C !B A)+(!D C B !A)+(!D C B A)), LSE_LINE_FILE_ID=3, LSE_LCOL=13, LSE_RCOL=44, LSE_LLINE=32, LSE_RLINE=32 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(11[2:53])
    defparam I1.init = 16'b0000000011111111;
    
endmodule
//
// Verilog Description of module inverter_U142
//

module inverter_U142 (\notGate[870]_keep , \notGate[871] ) /* synthesis syn_module_defined=1 */ ;
    input \notGate[870]_keep ;
    output \notGate[871] ;
    
    wire \notGate[870]_keep  /* synthesis alspreserve=1 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(25[15:22])
    
    LUT4 I1 (.A(\notGate[870]_keep ), .B(\notGate[870]_keep ), .C(\notGate[870]_keep ), 
         .D(\notGate[870]_keep ), .Z(\notGate[871] )) /* synthesis syn_instantiated=1, lut_function=((!D !C !B !A)+(!D !C !B A)+(!D !C B !A)+(!D !C B A)+(!D C !B !A)+(!D C !B A)+(!D C B !A)+(!D C B A)), LSE_LINE_FILE_ID=3, LSE_LCOL=13, LSE_RCOL=44, LSE_LLINE=32, LSE_RLINE=32 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(11[2:53])
    defparam I1.init = 16'b0000000011111111;
    
endmodule
//
// Verilog Description of module inverter_U143
//

module inverter_U143 (\notGate[869]_keep , \notGate[870] ) /* synthesis syn_module_defined=1 */ ;
    input \notGate[869]_keep ;
    output \notGate[870] ;
    
    wire \notGate[869]_keep  /* synthesis alspreserve=1 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(25[15:22])
    
    LUT4 I1 (.A(\notGate[869]_keep ), .B(\notGate[869]_keep ), .C(\notGate[869]_keep ), 
         .D(\notGate[869]_keep ), .Z(\notGate[870] )) /* synthesis syn_instantiated=1, lut_function=((!D !C !B !A)+(!D !C !B A)+(!D !C B !A)+(!D !C B A)+(!D C !B !A)+(!D C !B A)+(!D C B !A)+(!D C B A)), LSE_LINE_FILE_ID=3, LSE_LCOL=13, LSE_RCOL=44, LSE_LLINE=32, LSE_RLINE=32 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(11[2:53])
    defparam I1.init = 16'b0000000011111111;
    
endmodule
//
// Verilog Description of module inverter_U144
//

module inverter_U144 (\notGate[85]_keep , \notGate[86] ) /* synthesis syn_module_defined=1 */ ;
    input \notGate[85]_keep ;
    output \notGate[86] ;
    
    wire \notGate[85]_keep  /* synthesis alspreserve=1 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(25[15:22])
    
    LUT4 I1 (.A(\notGate[85]_keep ), .B(\notGate[85]_keep ), .C(\notGate[85]_keep ), 
         .D(\notGate[85]_keep ), .Z(\notGate[86] )) /* synthesis syn_instantiated=1, lut_function=((!D !C !B !A)+(!D !C !B A)+(!D !C B !A)+(!D !C B A)+(!D C !B !A)+(!D C !B A)+(!D C B !A)+(!D C B A)), LSE_LINE_FILE_ID=3, LSE_LCOL=13, LSE_RCOL=44, LSE_LLINE=32, LSE_RLINE=32 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(11[2:53])
    defparam I1.init = 16'b0000000011111111;
    
endmodule
//
// Verilog Description of module inverter_U145
//

module inverter_U145 (\notGate[868]_keep , \notGate[869] ) /* synthesis syn_module_defined=1 */ ;
    input \notGate[868]_keep ;
    output \notGate[869] ;
    
    wire \notGate[868]_keep  /* synthesis alspreserve=1 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(25[15:22])
    
    LUT4 I1 (.A(\notGate[868]_keep ), .B(\notGate[868]_keep ), .C(\notGate[868]_keep ), 
         .D(\notGate[868]_keep ), .Z(\notGate[869] )) /* synthesis syn_instantiated=1, lut_function=((!D !C !B !A)+(!D !C !B A)+(!D !C B !A)+(!D !C B A)+(!D C !B !A)+(!D C !B A)+(!D C B !A)+(!D C B A)), LSE_LINE_FILE_ID=3, LSE_LCOL=13, LSE_RCOL=44, LSE_LLINE=32, LSE_RLINE=32 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(11[2:53])
    defparam I1.init = 16'b0000000011111111;
    
endmodule
//
// Verilog Description of module inverter_U146
//

module inverter_U146 (\notGate[867]_keep , \notGate[868] ) /* synthesis syn_module_defined=1 */ ;
    input \notGate[867]_keep ;
    output \notGate[868] ;
    
    wire \notGate[867]_keep  /* synthesis alspreserve=1 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(25[15:22])
    
    LUT4 I1 (.A(\notGate[867]_keep ), .B(\notGate[867]_keep ), .C(\notGate[867]_keep ), 
         .D(\notGate[867]_keep ), .Z(\notGate[868] )) /* synthesis syn_instantiated=1, lut_function=((!D !C !B !A)+(!D !C !B A)+(!D !C B !A)+(!D !C B A)+(!D C !B !A)+(!D C !B A)+(!D C B !A)+(!D C B A)), LSE_LINE_FILE_ID=3, LSE_LCOL=13, LSE_RCOL=44, LSE_LLINE=32, LSE_RLINE=32 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(11[2:53])
    defparam I1.init = 16'b0000000011111111;
    
endmodule
//
// Verilog Description of module inverter_U147
//

module inverter_U147 (\notGate[866]_keep , \notGate[867] ) /* synthesis syn_module_defined=1 */ ;
    input \notGate[866]_keep ;
    output \notGate[867] ;
    
    wire \notGate[866]_keep  /* synthesis alspreserve=1 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(25[15:22])
    
    LUT4 I1 (.A(\notGate[866]_keep ), .B(\notGate[866]_keep ), .C(\notGate[866]_keep ), 
         .D(\notGate[866]_keep ), .Z(\notGate[867] )) /* synthesis syn_instantiated=1, lut_function=((!D !C !B !A)+(!D !C !B A)+(!D !C B !A)+(!D !C B A)+(!D C !B !A)+(!D C !B A)+(!D C B !A)+(!D C B A)), LSE_LINE_FILE_ID=3, LSE_LCOL=13, LSE_RCOL=44, LSE_LLINE=32, LSE_RLINE=32 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(11[2:53])
    defparam I1.init = 16'b0000000011111111;
    
endmodule
//
// Verilog Description of module inverter_U148
//

module inverter_U148 (\notGate[865]_keep , \notGate[866] ) /* synthesis syn_module_defined=1 */ ;
    input \notGate[865]_keep ;
    output \notGate[866] ;
    
    wire \notGate[865]_keep  /* synthesis alspreserve=1 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(25[15:22])
    
    LUT4 I1 (.A(\notGate[865]_keep ), .B(\notGate[865]_keep ), .C(\notGate[865]_keep ), 
         .D(\notGate[865]_keep ), .Z(\notGate[866] )) /* synthesis syn_instantiated=1, lut_function=((!D !C !B !A)+(!D !C !B A)+(!D !C B !A)+(!D !C B A)+(!D C !B !A)+(!D C !B A)+(!D C B !A)+(!D C B A)), LSE_LINE_FILE_ID=3, LSE_LCOL=13, LSE_RCOL=44, LSE_LLINE=32, LSE_RLINE=32 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(11[2:53])
    defparam I1.init = 16'b0000000011111111;
    
endmodule
//
// Verilog Description of module inverter_U149
//

module inverter_U149 (\notGate[864]_keep , \notGate[865] ) /* synthesis syn_module_defined=1 */ ;
    input \notGate[864]_keep ;
    output \notGate[865] ;
    
    wire \notGate[864]_keep  /* synthesis alspreserve=1 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(25[15:22])
    
    LUT4 I1 (.A(\notGate[864]_keep ), .B(\notGate[864]_keep ), .C(\notGate[864]_keep ), 
         .D(\notGate[864]_keep ), .Z(\notGate[865] )) /* synthesis syn_instantiated=1, lut_function=((!D !C !B !A)+(!D !C !B A)+(!D !C B !A)+(!D !C B A)+(!D C !B !A)+(!D C !B A)+(!D C B !A)+(!D C B A)), LSE_LINE_FILE_ID=3, LSE_LCOL=13, LSE_RCOL=44, LSE_LLINE=32, LSE_RLINE=32 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(11[2:53])
    defparam I1.init = 16'b0000000011111111;
    
endmodule
//
// Verilog Description of module inverter_U150
//

module inverter_U150 (\notGate[863]_keep , \notGate[864] ) /* synthesis syn_module_defined=1 */ ;
    input \notGate[863]_keep ;
    output \notGate[864] ;
    
    wire \notGate[863]_keep  /* synthesis alspreserve=1 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(25[15:22])
    
    LUT4 I1 (.A(\notGate[863]_keep ), .B(\notGate[863]_keep ), .C(\notGate[863]_keep ), 
         .D(\notGate[863]_keep ), .Z(\notGate[864] )) /* synthesis syn_instantiated=1, lut_function=((!D !C !B !A)+(!D !C !B A)+(!D !C B !A)+(!D !C B A)+(!D C !B !A)+(!D C !B A)+(!D C B !A)+(!D C B A)), LSE_LINE_FILE_ID=3, LSE_LCOL=13, LSE_RCOL=44, LSE_LLINE=32, LSE_RLINE=32 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(11[2:53])
    defparam I1.init = 16'b0000000011111111;
    
endmodule
//
// Verilog Description of module inverter_U151
//

module inverter_U151 (\notGate[862]_keep , \notGate[863] ) /* synthesis syn_module_defined=1 */ ;
    input \notGate[862]_keep ;
    output \notGate[863] ;
    
    wire \notGate[862]_keep  /* synthesis alspreserve=1 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(25[15:22])
    
    LUT4 I1 (.A(\notGate[862]_keep ), .B(\notGate[862]_keep ), .C(\notGate[862]_keep ), 
         .D(\notGate[862]_keep ), .Z(\notGate[863] )) /* synthesis syn_instantiated=1, lut_function=((!D !C !B !A)+(!D !C !B A)+(!D !C B !A)+(!D !C B A)+(!D C !B !A)+(!D C !B A)+(!D C B !A)+(!D C B A)), LSE_LINE_FILE_ID=3, LSE_LCOL=13, LSE_RCOL=44, LSE_LLINE=32, LSE_RLINE=32 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(11[2:53])
    defparam I1.init = 16'b0000000011111111;
    
endmodule
//
// Verilog Description of module inverter_U152
//

module inverter_U152 (\notGate[861]_keep , \notGate[862] ) /* synthesis syn_module_defined=1 */ ;
    input \notGate[861]_keep ;
    output \notGate[862] ;
    
    wire \notGate[861]_keep  /* synthesis alspreserve=1 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(25[15:22])
    
    LUT4 I1 (.A(\notGate[861]_keep ), .B(\notGate[861]_keep ), .C(\notGate[861]_keep ), 
         .D(\notGate[861]_keep ), .Z(\notGate[862] )) /* synthesis syn_instantiated=1, lut_function=((!D !C !B !A)+(!D !C !B A)+(!D !C B !A)+(!D !C B A)+(!D C !B !A)+(!D C !B A)+(!D C B !A)+(!D C B A)), LSE_LINE_FILE_ID=3, LSE_LCOL=13, LSE_RCOL=44, LSE_LLINE=32, LSE_RLINE=32 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(11[2:53])
    defparam I1.init = 16'b0000000011111111;
    
endmodule
//
// Verilog Description of module inverter_U153
//

module inverter_U153 (\notGate[860]_keep , \notGate[861] ) /* synthesis syn_module_defined=1 */ ;
    input \notGate[860]_keep ;
    output \notGate[861] ;
    
    wire \notGate[860]_keep  /* synthesis alspreserve=1 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(25[15:22])
    
    LUT4 I1 (.A(\notGate[860]_keep ), .B(\notGate[860]_keep ), .C(\notGate[860]_keep ), 
         .D(\notGate[860]_keep ), .Z(\notGate[861] )) /* synthesis syn_instantiated=1, lut_function=((!D !C !B !A)+(!D !C !B A)+(!D !C B !A)+(!D !C B A)+(!D C !B !A)+(!D C !B A)+(!D C B !A)+(!D C B A)), LSE_LINE_FILE_ID=3, LSE_LCOL=13, LSE_RCOL=44, LSE_LLINE=32, LSE_RLINE=32 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(11[2:53])
    defparam I1.init = 16'b0000000011111111;
    
endmodule
//
// Verilog Description of module inverter_U154
//

module inverter_U154 (\notGate[859]_keep , \notGate[860] ) /* synthesis syn_module_defined=1 */ ;
    input \notGate[859]_keep ;
    output \notGate[860] ;
    
    wire \notGate[859]_keep  /* synthesis alspreserve=1 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(25[15:22])
    
    LUT4 I1 (.A(\notGate[859]_keep ), .B(\notGate[859]_keep ), .C(\notGate[859]_keep ), 
         .D(\notGate[859]_keep ), .Z(\notGate[860] )) /* synthesis syn_instantiated=1, lut_function=((!D !C !B !A)+(!D !C !B A)+(!D !C B !A)+(!D !C B A)+(!D C !B !A)+(!D C !B A)+(!D C B !A)+(!D C B A)), LSE_LINE_FILE_ID=3, LSE_LCOL=13, LSE_RCOL=44, LSE_LLINE=32, LSE_RLINE=32 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(11[2:53])
    defparam I1.init = 16'b0000000011111111;
    
endmodule
//
// Verilog Description of module inverter_U155
//

module inverter_U155 (\notGate[84]_keep , \notGate[85] ) /* synthesis syn_module_defined=1 */ ;
    input \notGate[84]_keep ;
    output \notGate[85] ;
    
    wire \notGate[84]_keep  /* synthesis alspreserve=1 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(25[15:22])
    
    LUT4 I1 (.A(\notGate[84]_keep ), .B(\notGate[84]_keep ), .C(\notGate[84]_keep ), 
         .D(\notGate[84]_keep ), .Z(\notGate[85] )) /* synthesis syn_instantiated=1, lut_function=((!D !C !B !A)+(!D !C !B A)+(!D !C B !A)+(!D !C B A)+(!D C !B !A)+(!D C !B A)+(!D C B !A)+(!D C B A)), LSE_LINE_FILE_ID=3, LSE_LCOL=13, LSE_RCOL=44, LSE_LLINE=32, LSE_RLINE=32 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(11[2:53])
    defparam I1.init = 16'b0000000011111111;
    
endmodule
//
// Verilog Description of module inverter_U156
//

module inverter_U156 (\notGate[858]_keep , \notGate[859] ) /* synthesis syn_module_defined=1 */ ;
    input \notGate[858]_keep ;
    output \notGate[859] ;
    
    wire \notGate[858]_keep  /* synthesis alspreserve=1 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(25[15:22])
    
    LUT4 I1 (.A(\notGate[858]_keep ), .B(\notGate[858]_keep ), .C(\notGate[858]_keep ), 
         .D(\notGate[858]_keep ), .Z(\notGate[859] )) /* synthesis syn_instantiated=1, lut_function=((!D !C !B !A)+(!D !C !B A)+(!D !C B !A)+(!D !C B A)+(!D C !B !A)+(!D C !B A)+(!D C B !A)+(!D C B A)), LSE_LINE_FILE_ID=3, LSE_LCOL=13, LSE_RCOL=44, LSE_LLINE=32, LSE_RLINE=32 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(11[2:53])
    defparam I1.init = 16'b0000000011111111;
    
endmodule
//
// Verilog Description of module inverter_U157
//

module inverter_U157 (\notGate[857]_keep , \notGate[858] ) /* synthesis syn_module_defined=1 */ ;
    input \notGate[857]_keep ;
    output \notGate[858] ;
    
    wire \notGate[857]_keep  /* synthesis alspreserve=1 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(25[15:22])
    
    LUT4 I1 (.A(\notGate[857]_keep ), .B(\notGate[857]_keep ), .C(\notGate[857]_keep ), 
         .D(\notGate[857]_keep ), .Z(\notGate[858] )) /* synthesis syn_instantiated=1, lut_function=((!D !C !B !A)+(!D !C !B A)+(!D !C B !A)+(!D !C B A)+(!D C !B !A)+(!D C !B A)+(!D C B !A)+(!D C B A)), LSE_LINE_FILE_ID=3, LSE_LCOL=13, LSE_RCOL=44, LSE_LLINE=32, LSE_RLINE=32 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(11[2:53])
    defparam I1.init = 16'b0000000011111111;
    
endmodule
//
// Verilog Description of module inverter_U158
//

module inverter_U158 (\notGate[856]_keep , \notGate[857] ) /* synthesis syn_module_defined=1 */ ;
    input \notGate[856]_keep ;
    output \notGate[857] ;
    
    wire \notGate[856]_keep  /* synthesis alspreserve=1 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(25[15:22])
    
    LUT4 I1 (.A(\notGate[856]_keep ), .B(\notGate[856]_keep ), .C(\notGate[856]_keep ), 
         .D(\notGate[856]_keep ), .Z(\notGate[857] )) /* synthesis syn_instantiated=1, lut_function=((!D !C !B !A)+(!D !C !B A)+(!D !C B !A)+(!D !C B A)+(!D C !B !A)+(!D C !B A)+(!D C B !A)+(!D C B A)), LSE_LINE_FILE_ID=3, LSE_LCOL=13, LSE_RCOL=44, LSE_LLINE=32, LSE_RLINE=32 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(11[2:53])
    defparam I1.init = 16'b0000000011111111;
    
endmodule
//
// Verilog Description of module inverter_U159
//

module inverter_U159 (\notGate[855]_keep , \notGate[856] ) /* synthesis syn_module_defined=1 */ ;
    input \notGate[855]_keep ;
    output \notGate[856] ;
    
    wire \notGate[855]_keep  /* synthesis alspreserve=1 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(25[15:22])
    
    LUT4 I1 (.A(\notGate[855]_keep ), .B(\notGate[855]_keep ), .C(\notGate[855]_keep ), 
         .D(\notGate[855]_keep ), .Z(\notGate[856] )) /* synthesis syn_instantiated=1, lut_function=((!D !C !B !A)+(!D !C !B A)+(!D !C B !A)+(!D !C B A)+(!D C !B !A)+(!D C !B A)+(!D C B !A)+(!D C B A)), LSE_LINE_FILE_ID=3, LSE_LCOL=13, LSE_RCOL=44, LSE_LLINE=32, LSE_RLINE=32 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(11[2:53])
    defparam I1.init = 16'b0000000011111111;
    
endmodule
//
// Verilog Description of module inverter_U160
//

module inverter_U160 (\notGate[854]_keep , \notGate[855] ) /* synthesis syn_module_defined=1 */ ;
    input \notGate[854]_keep ;
    output \notGate[855] ;
    
    wire \notGate[854]_keep  /* synthesis alspreserve=1 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(25[15:22])
    
    LUT4 I1 (.A(\notGate[854]_keep ), .B(\notGate[854]_keep ), .C(\notGate[854]_keep ), 
         .D(\notGate[854]_keep ), .Z(\notGate[855] )) /* synthesis syn_instantiated=1, lut_function=((!D !C !B !A)+(!D !C !B A)+(!D !C B !A)+(!D !C B A)+(!D C !B !A)+(!D C !B A)+(!D C B !A)+(!D C B A)), LSE_LINE_FILE_ID=3, LSE_LCOL=13, LSE_RCOL=44, LSE_LLINE=32, LSE_RLINE=32 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(11[2:53])
    defparam I1.init = 16'b0000000011111111;
    
endmodule
//
// Verilog Description of module inverter_U161
//

module inverter_U161 (\notGate[853]_keep , \notGate[854] ) /* synthesis syn_module_defined=1 */ ;
    input \notGate[853]_keep ;
    output \notGate[854] ;
    
    wire \notGate[853]_keep  /* synthesis alspreserve=1 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(25[15:22])
    
    LUT4 I1 (.A(\notGate[853]_keep ), .B(\notGate[853]_keep ), .C(\notGate[853]_keep ), 
         .D(\notGate[853]_keep ), .Z(\notGate[854] )) /* synthesis syn_instantiated=1, lut_function=((!D !C !B !A)+(!D !C !B A)+(!D !C B !A)+(!D !C B A)+(!D C !B !A)+(!D C !B A)+(!D C B !A)+(!D C B A)), LSE_LINE_FILE_ID=3, LSE_LCOL=13, LSE_RCOL=44, LSE_LLINE=32, LSE_RLINE=32 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(11[2:53])
    defparam I1.init = 16'b0000000011111111;
    
endmodule
//
// Verilog Description of module inverter_U162
//

module inverter_U162 (\notGate[852]_keep , \notGate[853] ) /* synthesis syn_module_defined=1 */ ;
    input \notGate[852]_keep ;
    output \notGate[853] ;
    
    wire \notGate[852]_keep  /* synthesis alspreserve=1 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(25[15:22])
    
    LUT4 I1 (.A(\notGate[852]_keep ), .B(\notGate[852]_keep ), .C(\notGate[852]_keep ), 
         .D(\notGate[852]_keep ), .Z(\notGate[853] )) /* synthesis syn_instantiated=1, lut_function=((!D !C !B !A)+(!D !C !B A)+(!D !C B !A)+(!D !C B A)+(!D C !B !A)+(!D C !B A)+(!D C B !A)+(!D C B A)), LSE_LINE_FILE_ID=3, LSE_LCOL=13, LSE_RCOL=44, LSE_LLINE=32, LSE_RLINE=32 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(11[2:53])
    defparam I1.init = 16'b0000000011111111;
    
endmodule
//
// Verilog Description of module inverter_U163
//

module inverter_U163 (\notGate[851]_keep , \notGate[852] ) /* synthesis syn_module_defined=1 */ ;
    input \notGate[851]_keep ;
    output \notGate[852] ;
    
    wire \notGate[851]_keep  /* synthesis alspreserve=1 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(25[15:22])
    
    LUT4 I1 (.A(\notGate[851]_keep ), .B(\notGate[851]_keep ), .C(\notGate[851]_keep ), 
         .D(\notGate[851]_keep ), .Z(\notGate[852] )) /* synthesis syn_instantiated=1, lut_function=((!D !C !B !A)+(!D !C !B A)+(!D !C B !A)+(!D !C B A)+(!D C !B !A)+(!D C !B A)+(!D C B !A)+(!D C B A)), LSE_LINE_FILE_ID=3, LSE_LCOL=13, LSE_RCOL=44, LSE_LLINE=32, LSE_RLINE=32 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(11[2:53])
    defparam I1.init = 16'b0000000011111111;
    
endmodule
//
// Verilog Description of module inverter_U164
//

module inverter_U164 (\notGate[850]_keep , \notGate[851] ) /* synthesis syn_module_defined=1 */ ;
    input \notGate[850]_keep ;
    output \notGate[851] ;
    
    wire \notGate[850]_keep  /* synthesis alspreserve=1 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(25[15:22])
    
    LUT4 I1 (.A(\notGate[850]_keep ), .B(\notGate[850]_keep ), .C(\notGate[850]_keep ), 
         .D(\notGate[850]_keep ), .Z(\notGate[851] )) /* synthesis syn_instantiated=1, lut_function=((!D !C !B !A)+(!D !C !B A)+(!D !C B !A)+(!D !C B A)+(!D C !B !A)+(!D C !B A)+(!D C B !A)+(!D C B A)), LSE_LINE_FILE_ID=3, LSE_LCOL=13, LSE_RCOL=44, LSE_LLINE=32, LSE_RLINE=32 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(11[2:53])
    defparam I1.init = 16'b0000000011111111;
    
endmodule
//
// Verilog Description of module inverter_U165
//

module inverter_U165 (\notGate[849]_keep , \notGate[850] ) /* synthesis syn_module_defined=1 */ ;
    input \notGate[849]_keep ;
    output \notGate[850] ;
    
    wire \notGate[849]_keep  /* synthesis alspreserve=1 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(25[15:22])
    
    LUT4 I1 (.A(\notGate[849]_keep ), .B(\notGate[849]_keep ), .C(\notGate[849]_keep ), 
         .D(\notGate[849]_keep ), .Z(\notGate[850] )) /* synthesis syn_instantiated=1, lut_function=((!D !C !B !A)+(!D !C !B A)+(!D !C B !A)+(!D !C B A)+(!D C !B !A)+(!D C !B A)+(!D C B !A)+(!D C B A)), LSE_LINE_FILE_ID=3, LSE_LCOL=13, LSE_RCOL=44, LSE_LLINE=32, LSE_RLINE=32 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(11[2:53])
    defparam I1.init = 16'b0000000011111111;
    
endmodule
//
// Verilog Description of module inverter_U166
//

module inverter_U166 (\notGate[83]_keep , \notGate[84] ) /* synthesis syn_module_defined=1 */ ;
    input \notGate[83]_keep ;
    output \notGate[84] ;
    
    wire \notGate[83]_keep  /* synthesis alspreserve=1 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(25[15:22])
    
    LUT4 I1 (.A(\notGate[83]_keep ), .B(\notGate[83]_keep ), .C(\notGate[83]_keep ), 
         .D(\notGate[83]_keep ), .Z(\notGate[84] )) /* synthesis syn_instantiated=1, lut_function=((!D !C !B !A)+(!D !C !B A)+(!D !C B !A)+(!D !C B A)+(!D C !B !A)+(!D C !B A)+(!D C B !A)+(!D C B A)), LSE_LINE_FILE_ID=3, LSE_LCOL=13, LSE_RCOL=44, LSE_LLINE=32, LSE_RLINE=32 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(11[2:53])
    defparam I1.init = 16'b0000000011111111;
    
endmodule
//
// Verilog Description of module inverter_U167
//

module inverter_U167 (\notGate[848]_keep , \notGate[849] ) /* synthesis syn_module_defined=1 */ ;
    input \notGate[848]_keep ;
    output \notGate[849] ;
    
    wire \notGate[848]_keep  /* synthesis alspreserve=1 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(25[15:22])
    
    LUT4 I1 (.A(\notGate[848]_keep ), .B(\notGate[848]_keep ), .C(\notGate[848]_keep ), 
         .D(\notGate[848]_keep ), .Z(\notGate[849] )) /* synthesis syn_instantiated=1, lut_function=((!D !C !B !A)+(!D !C !B A)+(!D !C B !A)+(!D !C B A)+(!D C !B !A)+(!D C !B A)+(!D C B !A)+(!D C B A)), LSE_LINE_FILE_ID=3, LSE_LCOL=13, LSE_RCOL=44, LSE_LLINE=32, LSE_RLINE=32 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(11[2:53])
    defparam I1.init = 16'b0000000011111111;
    
endmodule
//
// Verilog Description of module inverter_U168
//

module inverter_U168 (\notGate[847]_keep , \notGate[848] ) /* synthesis syn_module_defined=1 */ ;
    input \notGate[847]_keep ;
    output \notGate[848] ;
    
    wire \notGate[847]_keep  /* synthesis alspreserve=1 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(25[15:22])
    
    LUT4 I1 (.A(\notGate[847]_keep ), .B(\notGate[847]_keep ), .C(\notGate[847]_keep ), 
         .D(\notGate[847]_keep ), .Z(\notGate[848] )) /* synthesis syn_instantiated=1, lut_function=((!D !C !B !A)+(!D !C !B A)+(!D !C B !A)+(!D !C B A)+(!D C !B !A)+(!D C !B A)+(!D C B !A)+(!D C B A)), LSE_LINE_FILE_ID=3, LSE_LCOL=13, LSE_RCOL=44, LSE_LLINE=32, LSE_RLINE=32 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(11[2:53])
    defparam I1.init = 16'b0000000011111111;
    
endmodule
//
// Verilog Description of module inverter_U169
//

module inverter_U169 (\notGate[846]_keep , \notGate[847] ) /* synthesis syn_module_defined=1 */ ;
    input \notGate[846]_keep ;
    output \notGate[847] ;
    
    wire \notGate[846]_keep  /* synthesis alspreserve=1 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(25[15:22])
    
    LUT4 I1 (.A(\notGate[846]_keep ), .B(\notGate[846]_keep ), .C(\notGate[846]_keep ), 
         .D(\notGate[846]_keep ), .Z(\notGate[847] )) /* synthesis syn_instantiated=1, lut_function=((!D !C !B !A)+(!D !C !B A)+(!D !C B !A)+(!D !C B A)+(!D C !B !A)+(!D C !B A)+(!D C B !A)+(!D C B A)), LSE_LINE_FILE_ID=3, LSE_LCOL=13, LSE_RCOL=44, LSE_LLINE=32, LSE_RLINE=32 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(11[2:53])
    defparam I1.init = 16'b0000000011111111;
    
endmodule
//
// Verilog Description of module inverter_U170
//

module inverter_U170 (\notGate[845]_keep , \notGate[846] ) /* synthesis syn_module_defined=1 */ ;
    input \notGate[845]_keep ;
    output \notGate[846] ;
    
    wire \notGate[845]_keep  /* synthesis alspreserve=1 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(25[15:22])
    
    LUT4 I1 (.A(\notGate[845]_keep ), .B(\notGate[845]_keep ), .C(\notGate[845]_keep ), 
         .D(\notGate[845]_keep ), .Z(\notGate[846] )) /* synthesis syn_instantiated=1, lut_function=((!D !C !B !A)+(!D !C !B A)+(!D !C B !A)+(!D !C B A)+(!D C !B !A)+(!D C !B A)+(!D C B !A)+(!D C B A)), LSE_LINE_FILE_ID=3, LSE_LCOL=13, LSE_RCOL=44, LSE_LLINE=32, LSE_RLINE=32 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(11[2:53])
    defparam I1.init = 16'b0000000011111111;
    
endmodule
//
// Verilog Description of module inverter_U171
//

module inverter_U171 (\notGate[844]_keep , \notGate[845] ) /* synthesis syn_module_defined=1 */ ;
    input \notGate[844]_keep ;
    output \notGate[845] ;
    
    wire \notGate[844]_keep  /* synthesis alspreserve=1 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(25[15:22])
    
    LUT4 I1 (.A(\notGate[844]_keep ), .B(\notGate[844]_keep ), .C(\notGate[844]_keep ), 
         .D(\notGate[844]_keep ), .Z(\notGate[845] )) /* synthesis syn_instantiated=1, lut_function=((!D !C !B !A)+(!D !C !B A)+(!D !C B !A)+(!D !C B A)+(!D C !B !A)+(!D C !B A)+(!D C B !A)+(!D C B A)), LSE_LINE_FILE_ID=3, LSE_LCOL=13, LSE_RCOL=44, LSE_LLINE=32, LSE_RLINE=32 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(11[2:53])
    defparam I1.init = 16'b0000000011111111;
    
endmodule
//
// Verilog Description of module inverter_U172
//

module inverter_U172 (\notGate[843]_keep , \notGate[844] ) /* synthesis syn_module_defined=1 */ ;
    input \notGate[843]_keep ;
    output \notGate[844] ;
    
    wire \notGate[843]_keep  /* synthesis alspreserve=1 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(25[15:22])
    
    LUT4 I1 (.A(\notGate[843]_keep ), .B(\notGate[843]_keep ), .C(\notGate[843]_keep ), 
         .D(\notGate[843]_keep ), .Z(\notGate[844] )) /* synthesis syn_instantiated=1, lut_function=((!D !C !B !A)+(!D !C !B A)+(!D !C B !A)+(!D !C B A)+(!D C !B !A)+(!D C !B A)+(!D C B !A)+(!D C B A)), LSE_LINE_FILE_ID=3, LSE_LCOL=13, LSE_RCOL=44, LSE_LLINE=32, LSE_RLINE=32 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(11[2:53])
    defparam I1.init = 16'b0000000011111111;
    
endmodule
//
// Verilog Description of module inverter_U173
//

module inverter_U173 (\notGate[842]_keep , \notGate[843] ) /* synthesis syn_module_defined=1 */ ;
    input \notGate[842]_keep ;
    output \notGate[843] ;
    
    wire \notGate[842]_keep  /* synthesis alspreserve=1 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(25[15:22])
    
    LUT4 I1 (.A(\notGate[842]_keep ), .B(\notGate[842]_keep ), .C(\notGate[842]_keep ), 
         .D(\notGate[842]_keep ), .Z(\notGate[843] )) /* synthesis syn_instantiated=1, lut_function=((!D !C !B !A)+(!D !C !B A)+(!D !C B !A)+(!D !C B A)+(!D C !B !A)+(!D C !B A)+(!D C B !A)+(!D C B A)), LSE_LINE_FILE_ID=3, LSE_LCOL=13, LSE_RCOL=44, LSE_LLINE=32, LSE_RLINE=32 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(11[2:53])
    defparam I1.init = 16'b0000000011111111;
    
endmodule
//
// Verilog Description of module inverter_U174
//

module inverter_U174 (\notGate[841]_keep , \notGate[842] ) /* synthesis syn_module_defined=1 */ ;
    input \notGate[841]_keep ;
    output \notGate[842] ;
    
    wire \notGate[841]_keep  /* synthesis alspreserve=1 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(25[15:22])
    
    LUT4 I1 (.A(\notGate[841]_keep ), .B(\notGate[841]_keep ), .C(\notGate[841]_keep ), 
         .D(\notGate[841]_keep ), .Z(\notGate[842] )) /* synthesis syn_instantiated=1, lut_function=((!D !C !B !A)+(!D !C !B A)+(!D !C B !A)+(!D !C B A)+(!D C !B !A)+(!D C !B A)+(!D C B !A)+(!D C B A)), LSE_LINE_FILE_ID=3, LSE_LCOL=13, LSE_RCOL=44, LSE_LLINE=32, LSE_RLINE=32 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(11[2:53])
    defparam I1.init = 16'b0000000011111111;
    
endmodule
//
// Verilog Description of module inverter_U175
//

module inverter_U175 (\notGate[840]_keep , \notGate[841] ) /* synthesis syn_module_defined=1 */ ;
    input \notGate[840]_keep ;
    output \notGate[841] ;
    
    wire \notGate[840]_keep  /* synthesis alspreserve=1 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(25[15:22])
    
    LUT4 I1 (.A(\notGate[840]_keep ), .B(\notGate[840]_keep ), .C(\notGate[840]_keep ), 
         .D(\notGate[840]_keep ), .Z(\notGate[841] )) /* synthesis syn_instantiated=1, lut_function=((!D !C !B !A)+(!D !C !B A)+(!D !C B !A)+(!D !C B A)+(!D C !B !A)+(!D C !B A)+(!D C B !A)+(!D C B A)), LSE_LINE_FILE_ID=3, LSE_LCOL=13, LSE_RCOL=44, LSE_LLINE=32, LSE_RLINE=32 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(11[2:53])
    defparam I1.init = 16'b0000000011111111;
    
endmodule
//
// Verilog Description of module inverter_U176
//

module inverter_U176 (\notGate[839]_keep , \notGate[840] ) /* synthesis syn_module_defined=1 */ ;
    input \notGate[839]_keep ;
    output \notGate[840] ;
    
    wire \notGate[839]_keep  /* synthesis alspreserve=1 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(25[15:22])
    
    LUT4 I1 (.A(\notGate[839]_keep ), .B(\notGate[839]_keep ), .C(\notGate[839]_keep ), 
         .D(\notGate[839]_keep ), .Z(\notGate[840] )) /* synthesis syn_instantiated=1, lut_function=((!D !C !B !A)+(!D !C !B A)+(!D !C B !A)+(!D !C B A)+(!D C !B !A)+(!D C !B A)+(!D C B !A)+(!D C B A)), LSE_LINE_FILE_ID=3, LSE_LCOL=13, LSE_RCOL=44, LSE_LLINE=32, LSE_RLINE=32 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(11[2:53])
    defparam I1.init = 16'b0000000011111111;
    
endmodule
//
// Verilog Description of module inverter_U177
//

module inverter_U177 (\notGate[82]_keep , \notGate[83] ) /* synthesis syn_module_defined=1 */ ;
    input \notGate[82]_keep ;
    output \notGate[83] ;
    
    wire \notGate[82]_keep  /* synthesis alspreserve=1 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(25[15:22])
    
    LUT4 I1 (.A(\notGate[82]_keep ), .B(\notGate[82]_keep ), .C(\notGate[82]_keep ), 
         .D(\notGate[82]_keep ), .Z(\notGate[83] )) /* synthesis syn_instantiated=1, lut_function=((!D !C !B !A)+(!D !C !B A)+(!D !C B !A)+(!D !C B A)+(!D C !B !A)+(!D C !B A)+(!D C B !A)+(!D C B A)), LSE_LINE_FILE_ID=3, LSE_LCOL=13, LSE_RCOL=44, LSE_LLINE=32, LSE_RLINE=32 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(11[2:53])
    defparam I1.init = 16'b0000000011111111;
    
endmodule
//
// Verilog Description of module inverter_U178
//

module inverter_U178 (\notGate[838]_keep , \notGate[839] ) /* synthesis syn_module_defined=1 */ ;
    input \notGate[838]_keep ;
    output \notGate[839] ;
    
    wire \notGate[838]_keep  /* synthesis alspreserve=1 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(25[15:22])
    
    LUT4 I1 (.A(\notGate[838]_keep ), .B(\notGate[838]_keep ), .C(\notGate[838]_keep ), 
         .D(\notGate[838]_keep ), .Z(\notGate[839] )) /* synthesis syn_instantiated=1, lut_function=((!D !C !B !A)+(!D !C !B A)+(!D !C B !A)+(!D !C B A)+(!D C !B !A)+(!D C !B A)+(!D C B !A)+(!D C B A)), LSE_LINE_FILE_ID=3, LSE_LCOL=13, LSE_RCOL=44, LSE_LLINE=32, LSE_RLINE=32 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(11[2:53])
    defparam I1.init = 16'b0000000011111111;
    
endmodule
//
// Verilog Description of module inverter_U179
//

module inverter_U179 (\notGate[837]_keep , \notGate[838] ) /* synthesis syn_module_defined=1 */ ;
    input \notGate[837]_keep ;
    output \notGate[838] ;
    
    wire \notGate[837]_keep  /* synthesis alspreserve=1 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(25[15:22])
    
    LUT4 I1 (.A(\notGate[837]_keep ), .B(\notGate[837]_keep ), .C(\notGate[837]_keep ), 
         .D(\notGate[837]_keep ), .Z(\notGate[838] )) /* synthesis syn_instantiated=1, lut_function=((!D !C !B !A)+(!D !C !B A)+(!D !C B !A)+(!D !C B A)+(!D C !B !A)+(!D C !B A)+(!D C B !A)+(!D C B A)), LSE_LINE_FILE_ID=3, LSE_LCOL=13, LSE_RCOL=44, LSE_LLINE=32, LSE_RLINE=32 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(11[2:53])
    defparam I1.init = 16'b0000000011111111;
    
endmodule
//
// Verilog Description of module inverter_U180
//

module inverter_U180 (\notGate[836]_keep , \notGate[837] ) /* synthesis syn_module_defined=1 */ ;
    input \notGate[836]_keep ;
    output \notGate[837] ;
    
    wire \notGate[836]_keep  /* synthesis alspreserve=1 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(25[15:22])
    
    LUT4 I1 (.A(\notGate[836]_keep ), .B(\notGate[836]_keep ), .C(\notGate[836]_keep ), 
         .D(\notGate[836]_keep ), .Z(\notGate[837] )) /* synthesis syn_instantiated=1, lut_function=((!D !C !B !A)+(!D !C !B A)+(!D !C B !A)+(!D !C B A)+(!D C !B !A)+(!D C !B A)+(!D C B !A)+(!D C B A)), LSE_LINE_FILE_ID=3, LSE_LCOL=13, LSE_RCOL=44, LSE_LLINE=32, LSE_RLINE=32 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(11[2:53])
    defparam I1.init = 16'b0000000011111111;
    
endmodule
//
// Verilog Description of module inverter_U181
//

module inverter_U181 (\notGate[835]_keep , \notGate[836] ) /* synthesis syn_module_defined=1 */ ;
    input \notGate[835]_keep ;
    output \notGate[836] ;
    
    wire \notGate[835]_keep  /* synthesis alspreserve=1 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(25[15:22])
    
    LUT4 I1 (.A(\notGate[835]_keep ), .B(\notGate[835]_keep ), .C(\notGate[835]_keep ), 
         .D(\notGate[835]_keep ), .Z(\notGate[836] )) /* synthesis syn_instantiated=1, lut_function=((!D !C !B !A)+(!D !C !B A)+(!D !C B !A)+(!D !C B A)+(!D C !B !A)+(!D C !B A)+(!D C B !A)+(!D C B A)), LSE_LINE_FILE_ID=3, LSE_LCOL=13, LSE_RCOL=44, LSE_LLINE=32, LSE_RLINE=32 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(11[2:53])
    defparam I1.init = 16'b0000000011111111;
    
endmodule
//
// Verilog Description of module inverter_U182
//

module inverter_U182 (\notGate[834]_keep , \notGate[835] ) /* synthesis syn_module_defined=1 */ ;
    input \notGate[834]_keep ;
    output \notGate[835] ;
    
    wire \notGate[834]_keep  /* synthesis alspreserve=1 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(25[15:22])
    
    LUT4 I1 (.A(\notGate[834]_keep ), .B(\notGate[834]_keep ), .C(\notGate[834]_keep ), 
         .D(\notGate[834]_keep ), .Z(\notGate[835] )) /* synthesis syn_instantiated=1, lut_function=((!D !C !B !A)+(!D !C !B A)+(!D !C B !A)+(!D !C B A)+(!D C !B !A)+(!D C !B A)+(!D C B !A)+(!D C B A)), LSE_LINE_FILE_ID=3, LSE_LCOL=13, LSE_RCOL=44, LSE_LLINE=32, LSE_RLINE=32 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(11[2:53])
    defparam I1.init = 16'b0000000011111111;
    
endmodule
//
// Verilog Description of module inverter_U183
//

module inverter_U183 (\notGate[833]_keep , \notGate[834] ) /* synthesis syn_module_defined=1 */ ;
    input \notGate[833]_keep ;
    output \notGate[834] ;
    
    wire \notGate[833]_keep  /* synthesis alspreserve=1 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(25[15:22])
    
    LUT4 I1 (.A(\notGate[833]_keep ), .B(\notGate[833]_keep ), .C(\notGate[833]_keep ), 
         .D(\notGate[833]_keep ), .Z(\notGate[834] )) /* synthesis syn_instantiated=1, lut_function=((!D !C !B !A)+(!D !C !B A)+(!D !C B !A)+(!D !C B A)+(!D C !B !A)+(!D C !B A)+(!D C B !A)+(!D C B A)), LSE_LINE_FILE_ID=3, LSE_LCOL=13, LSE_RCOL=44, LSE_LLINE=32, LSE_RLINE=32 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(11[2:53])
    defparam I1.init = 16'b0000000011111111;
    
endmodule
//
// Verilog Description of module inverter_U184
//

module inverter_U184 (\notGate[832]_keep , \notGate[833] ) /* synthesis syn_module_defined=1 */ ;
    input \notGate[832]_keep ;
    output \notGate[833] ;
    
    wire \notGate[832]_keep  /* synthesis alspreserve=1 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(25[15:22])
    
    LUT4 I1 (.A(\notGate[832]_keep ), .B(\notGate[832]_keep ), .C(\notGate[832]_keep ), 
         .D(\notGate[832]_keep ), .Z(\notGate[833] )) /* synthesis syn_instantiated=1, lut_function=((!D !C !B !A)+(!D !C !B A)+(!D !C B !A)+(!D !C B A)+(!D C !B !A)+(!D C !B A)+(!D C B !A)+(!D C B A)), LSE_LINE_FILE_ID=3, LSE_LCOL=13, LSE_RCOL=44, LSE_LLINE=32, LSE_RLINE=32 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(11[2:53])
    defparam I1.init = 16'b0000000011111111;
    
endmodule
//
// Verilog Description of module inverter_U185
//

module inverter_U185 (\notGate[831]_keep , \notGate[832] ) /* synthesis syn_module_defined=1 */ ;
    input \notGate[831]_keep ;
    output \notGate[832] ;
    
    wire \notGate[831]_keep  /* synthesis alspreserve=1 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(25[15:22])
    
    LUT4 I1 (.A(\notGate[831]_keep ), .B(\notGate[831]_keep ), .C(\notGate[831]_keep ), 
         .D(\notGate[831]_keep ), .Z(\notGate[832] )) /* synthesis syn_instantiated=1, lut_function=((!D !C !B !A)+(!D !C !B A)+(!D !C B !A)+(!D !C B A)+(!D C !B !A)+(!D C !B A)+(!D C B !A)+(!D C B A)), LSE_LINE_FILE_ID=3, LSE_LCOL=13, LSE_RCOL=44, LSE_LLINE=32, LSE_RLINE=32 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(11[2:53])
    defparam I1.init = 16'b0000000011111111;
    
endmodule
//
// Verilog Description of module inverter_U186
//

module inverter_U186 (\notGate[830]_keep , \notGate[831] ) /* synthesis syn_module_defined=1 */ ;
    input \notGate[830]_keep ;
    output \notGate[831] ;
    
    wire \notGate[830]_keep  /* synthesis alspreserve=1 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(25[15:22])
    
    LUT4 I1 (.A(\notGate[830]_keep ), .B(\notGate[830]_keep ), .C(\notGate[830]_keep ), 
         .D(\notGate[830]_keep ), .Z(\notGate[831] )) /* synthesis syn_instantiated=1, lut_function=((!D !C !B !A)+(!D !C !B A)+(!D !C B !A)+(!D !C B A)+(!D C !B !A)+(!D C !B A)+(!D C B !A)+(!D C B A)), LSE_LINE_FILE_ID=3, LSE_LCOL=13, LSE_RCOL=44, LSE_LLINE=32, LSE_RLINE=32 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(11[2:53])
    defparam I1.init = 16'b0000000011111111;
    
endmodule
//
// Verilog Description of module inverter_U187
//

module inverter_U187 (\notGate[829]_keep , \notGate[830] ) /* synthesis syn_module_defined=1 */ ;
    input \notGate[829]_keep ;
    output \notGate[830] ;
    
    wire \notGate[829]_keep  /* synthesis alspreserve=1 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(25[15:22])
    
    LUT4 I1 (.A(\notGate[829]_keep ), .B(\notGate[829]_keep ), .C(\notGate[829]_keep ), 
         .D(\notGate[829]_keep ), .Z(\notGate[830] )) /* synthesis syn_instantiated=1, lut_function=((!D !C !B !A)+(!D !C !B A)+(!D !C B !A)+(!D !C B A)+(!D C !B !A)+(!D C !B A)+(!D C B !A)+(!D C B A)), LSE_LINE_FILE_ID=3, LSE_LCOL=13, LSE_RCOL=44, LSE_LLINE=32, LSE_RLINE=32 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(11[2:53])
    defparam I1.init = 16'b0000000011111111;
    
endmodule
//
// Verilog Description of module inverter_U188
//

module inverter_U188 (\notGate[81]_keep , \notGate[82] ) /* synthesis syn_module_defined=1 */ ;
    input \notGate[81]_keep ;
    output \notGate[82] ;
    
    wire \notGate[81]_keep  /* synthesis alspreserve=1 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(25[15:22])
    
    LUT4 I1 (.A(\notGate[81]_keep ), .B(\notGate[81]_keep ), .C(\notGate[81]_keep ), 
         .D(\notGate[81]_keep ), .Z(\notGate[82] )) /* synthesis syn_instantiated=1, lut_function=((!D !C !B !A)+(!D !C !B A)+(!D !C B !A)+(!D !C B A)+(!D C !B !A)+(!D C !B A)+(!D C B !A)+(!D C B A)), LSE_LINE_FILE_ID=3, LSE_LCOL=13, LSE_RCOL=44, LSE_LLINE=32, LSE_RLINE=32 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(11[2:53])
    defparam I1.init = 16'b0000000011111111;
    
endmodule
//
// Verilog Description of module inverter_U189
//

module inverter_U189 (\notGate[828]_keep , \notGate[829] ) /* synthesis syn_module_defined=1 */ ;
    input \notGate[828]_keep ;
    output \notGate[829] ;
    
    wire \notGate[828]_keep  /* synthesis alspreserve=1 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(25[15:22])
    
    LUT4 I1 (.A(\notGate[828]_keep ), .B(\notGate[828]_keep ), .C(\notGate[828]_keep ), 
         .D(\notGate[828]_keep ), .Z(\notGate[829] )) /* synthesis syn_instantiated=1, lut_function=((!D !C !B !A)+(!D !C !B A)+(!D !C B !A)+(!D !C B A)+(!D C !B !A)+(!D C !B A)+(!D C B !A)+(!D C B A)), LSE_LINE_FILE_ID=3, LSE_LCOL=13, LSE_RCOL=44, LSE_LLINE=32, LSE_RLINE=32 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(11[2:53])
    defparam I1.init = 16'b0000000011111111;
    
endmodule
//
// Verilog Description of module inverter_U190
//

module inverter_U190 (\notGate[827]_keep , \notGate[828] ) /* synthesis syn_module_defined=1 */ ;
    input \notGate[827]_keep ;
    output \notGate[828] ;
    
    wire \notGate[827]_keep  /* synthesis alspreserve=1 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(25[15:22])
    
    LUT4 I1 (.A(\notGate[827]_keep ), .B(\notGate[827]_keep ), .C(\notGate[827]_keep ), 
         .D(\notGate[827]_keep ), .Z(\notGate[828] )) /* synthesis syn_instantiated=1, lut_function=((!D !C !B !A)+(!D !C !B A)+(!D !C B !A)+(!D !C B A)+(!D C !B !A)+(!D C !B A)+(!D C B !A)+(!D C B A)), LSE_LINE_FILE_ID=3, LSE_LCOL=13, LSE_RCOL=44, LSE_LLINE=32, LSE_RLINE=32 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(11[2:53])
    defparam I1.init = 16'b0000000011111111;
    
endmodule
//
// Verilog Description of module inverter_U191
//

module inverter_U191 (\notGate[826]_keep , \notGate[827] ) /* synthesis syn_module_defined=1 */ ;
    input \notGate[826]_keep ;
    output \notGate[827] ;
    
    wire \notGate[826]_keep  /* synthesis alspreserve=1 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(25[15:22])
    
    LUT4 I1 (.A(\notGate[826]_keep ), .B(\notGate[826]_keep ), .C(\notGate[826]_keep ), 
         .D(\notGate[826]_keep ), .Z(\notGate[827] )) /* synthesis syn_instantiated=1, lut_function=((!D !C !B !A)+(!D !C !B A)+(!D !C B !A)+(!D !C B A)+(!D C !B !A)+(!D C !B A)+(!D C B !A)+(!D C B A)), LSE_LINE_FILE_ID=3, LSE_LCOL=13, LSE_RCOL=44, LSE_LLINE=32, LSE_RLINE=32 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(11[2:53])
    defparam I1.init = 16'b0000000011111111;
    
endmodule
//
// Verilog Description of module inverter_U192
//

module inverter_U192 (\notGate[825]_keep , \notGate[826] ) /* synthesis syn_module_defined=1 */ ;
    input \notGate[825]_keep ;
    output \notGate[826] ;
    
    wire \notGate[825]_keep  /* synthesis alspreserve=1 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(25[15:22])
    
    LUT4 I1 (.A(\notGate[825]_keep ), .B(\notGate[825]_keep ), .C(\notGate[825]_keep ), 
         .D(\notGate[825]_keep ), .Z(\notGate[826] )) /* synthesis syn_instantiated=1, lut_function=((!D !C !B !A)+(!D !C !B A)+(!D !C B !A)+(!D !C B A)+(!D C !B !A)+(!D C !B A)+(!D C B !A)+(!D C B A)), LSE_LINE_FILE_ID=3, LSE_LCOL=13, LSE_RCOL=44, LSE_LLINE=32, LSE_RLINE=32 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(11[2:53])
    defparam I1.init = 16'b0000000011111111;
    
endmodule
//
// Verilog Description of module inverter_U193
//

module inverter_U193 (\notGate[824]_keep , \notGate[825] ) /* synthesis syn_module_defined=1 */ ;
    input \notGate[824]_keep ;
    output \notGate[825] ;
    
    wire \notGate[824]_keep  /* synthesis alspreserve=1 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(25[15:22])
    
    LUT4 I1 (.A(\notGate[824]_keep ), .B(\notGate[824]_keep ), .C(\notGate[824]_keep ), 
         .D(\notGate[824]_keep ), .Z(\notGate[825] )) /* synthesis syn_instantiated=1, lut_function=((!D !C !B !A)+(!D !C !B A)+(!D !C B !A)+(!D !C B A)+(!D C !B !A)+(!D C !B A)+(!D C B !A)+(!D C B A)), LSE_LINE_FILE_ID=3, LSE_LCOL=13, LSE_RCOL=44, LSE_LLINE=32, LSE_RLINE=32 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(11[2:53])
    defparam I1.init = 16'b0000000011111111;
    
endmodule
//
// Verilog Description of module inverter_U194
//

module inverter_U194 (\notGate[823]_keep , \notGate[824] ) /* synthesis syn_module_defined=1 */ ;
    input \notGate[823]_keep ;
    output \notGate[824] ;
    
    wire \notGate[823]_keep  /* synthesis alspreserve=1 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(25[15:22])
    
    LUT4 I1 (.A(\notGate[823]_keep ), .B(\notGate[823]_keep ), .C(\notGate[823]_keep ), 
         .D(\notGate[823]_keep ), .Z(\notGate[824] )) /* synthesis syn_instantiated=1, lut_function=((!D !C !B !A)+(!D !C !B A)+(!D !C B !A)+(!D !C B A)+(!D C !B !A)+(!D C !B A)+(!D C B !A)+(!D C B A)), LSE_LINE_FILE_ID=3, LSE_LCOL=13, LSE_RCOL=44, LSE_LLINE=32, LSE_RLINE=32 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(11[2:53])
    defparam I1.init = 16'b0000000011111111;
    
endmodule
//
// Verilog Description of module inverter_U195
//

module inverter_U195 (\notGate[822]_keep , \notGate[823] ) /* synthesis syn_module_defined=1 */ ;
    input \notGate[822]_keep ;
    output \notGate[823] ;
    
    wire \notGate[822]_keep  /* synthesis alspreserve=1 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(25[15:22])
    
    LUT4 I1 (.A(\notGate[822]_keep ), .B(\notGate[822]_keep ), .C(\notGate[822]_keep ), 
         .D(\notGate[822]_keep ), .Z(\notGate[823] )) /* synthesis syn_instantiated=1, lut_function=((!D !C !B !A)+(!D !C !B A)+(!D !C B !A)+(!D !C B A)+(!D C !B !A)+(!D C !B A)+(!D C B !A)+(!D C B A)), LSE_LINE_FILE_ID=3, LSE_LCOL=13, LSE_RCOL=44, LSE_LLINE=32, LSE_RLINE=32 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(11[2:53])
    defparam I1.init = 16'b0000000011111111;
    
endmodule
//
// Verilog Description of module inverter_U196
//

module inverter_U196 (\notGate[821]_keep , \notGate[822] ) /* synthesis syn_module_defined=1 */ ;
    input \notGate[821]_keep ;
    output \notGate[822] ;
    
    wire \notGate[821]_keep  /* synthesis alspreserve=1 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(25[15:22])
    
    LUT4 I1 (.A(\notGate[821]_keep ), .B(\notGate[821]_keep ), .C(\notGate[821]_keep ), 
         .D(\notGate[821]_keep ), .Z(\notGate[822] )) /* synthesis syn_instantiated=1, lut_function=((!D !C !B !A)+(!D !C !B A)+(!D !C B !A)+(!D !C B A)+(!D C !B !A)+(!D C !B A)+(!D C B !A)+(!D C B A)), LSE_LINE_FILE_ID=3, LSE_LCOL=13, LSE_RCOL=44, LSE_LLINE=32, LSE_RLINE=32 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(11[2:53])
    defparam I1.init = 16'b0000000011111111;
    
endmodule
//
// Verilog Description of module inverter_U197
//

module inverter_U197 (\notGate[820]_keep , \notGate[821] ) /* synthesis syn_module_defined=1 */ ;
    input \notGate[820]_keep ;
    output \notGate[821] ;
    
    wire \notGate[820]_keep  /* synthesis alspreserve=1 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(25[15:22])
    
    LUT4 I1 (.A(\notGate[820]_keep ), .B(\notGate[820]_keep ), .C(\notGate[820]_keep ), 
         .D(\notGate[820]_keep ), .Z(\notGate[821] )) /* synthesis syn_instantiated=1, lut_function=((!D !C !B !A)+(!D !C !B A)+(!D !C B !A)+(!D !C B A)+(!D C !B !A)+(!D C !B A)+(!D C B !A)+(!D C B A)), LSE_LINE_FILE_ID=3, LSE_LCOL=13, LSE_RCOL=44, LSE_LLINE=32, LSE_RLINE=32 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(11[2:53])
    defparam I1.init = 16'b0000000011111111;
    
endmodule
//
// Verilog Description of module inverter_U198
//

module inverter_U198 (\notGate[819]_keep , \notGate[820] ) /* synthesis syn_module_defined=1 */ ;
    input \notGate[819]_keep ;
    output \notGate[820] ;
    
    wire \notGate[819]_keep  /* synthesis alspreserve=1 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(25[15:22])
    
    LUT4 I1 (.A(\notGate[819]_keep ), .B(\notGate[819]_keep ), .C(\notGate[819]_keep ), 
         .D(\notGate[819]_keep ), .Z(\notGate[820] )) /* synthesis syn_instantiated=1, lut_function=((!D !C !B !A)+(!D !C !B A)+(!D !C B !A)+(!D !C B A)+(!D C !B !A)+(!D C !B A)+(!D C B !A)+(!D C B A)), LSE_LINE_FILE_ID=3, LSE_LCOL=13, LSE_RCOL=44, LSE_LLINE=32, LSE_RLINE=32 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(11[2:53])
    defparam I1.init = 16'b0000000011111111;
    
endmodule
//
// Verilog Description of module inverter_U199
//

module inverter_U199 (\notGate[80]_keep , \notGate[81] ) /* synthesis syn_module_defined=1 */ ;
    input \notGate[80]_keep ;
    output \notGate[81] ;
    
    wire \notGate[80]_keep  /* synthesis alspreserve=1 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(25[15:22])
    
    LUT4 I1 (.A(\notGate[80]_keep ), .B(\notGate[80]_keep ), .C(\notGate[80]_keep ), 
         .D(\notGate[80]_keep ), .Z(\notGate[81] )) /* synthesis syn_instantiated=1, lut_function=((!D !C !B !A)+(!D !C !B A)+(!D !C B !A)+(!D !C B A)+(!D C !B !A)+(!D C !B A)+(!D C B !A)+(!D C B A)), LSE_LINE_FILE_ID=3, LSE_LCOL=13, LSE_RCOL=44, LSE_LLINE=32, LSE_RLINE=32 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(11[2:53])
    defparam I1.init = 16'b0000000011111111;
    
endmodule
//
// Verilog Description of module inverter_U200
//

module inverter_U200 (\notGate[818]_keep , \notGate[819] ) /* synthesis syn_module_defined=1 */ ;
    input \notGate[818]_keep ;
    output \notGate[819] ;
    
    wire \notGate[818]_keep  /* synthesis alspreserve=1 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(25[15:22])
    
    LUT4 I1 (.A(\notGate[818]_keep ), .B(\notGate[818]_keep ), .C(\notGate[818]_keep ), 
         .D(\notGate[818]_keep ), .Z(\notGate[819] )) /* synthesis syn_instantiated=1, lut_function=((!D !C !B !A)+(!D !C !B A)+(!D !C B !A)+(!D !C B A)+(!D C !B !A)+(!D C !B A)+(!D C B !A)+(!D C B A)), LSE_LINE_FILE_ID=3, LSE_LCOL=13, LSE_RCOL=44, LSE_LLINE=32, LSE_RLINE=32 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(11[2:53])
    defparam I1.init = 16'b0000000011111111;
    
endmodule
//
// Verilog Description of module inverter_U201
//

module inverter_U201 (\notGate[817]_keep , \notGate[818] ) /* synthesis syn_module_defined=1 */ ;
    input \notGate[817]_keep ;
    output \notGate[818] ;
    
    wire \notGate[817]_keep  /* synthesis alspreserve=1 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(25[15:22])
    
    LUT4 I1 (.A(\notGate[817]_keep ), .B(\notGate[817]_keep ), .C(\notGate[817]_keep ), 
         .D(\notGate[817]_keep ), .Z(\notGate[818] )) /* synthesis syn_instantiated=1, lut_function=((!D !C !B !A)+(!D !C !B A)+(!D !C B !A)+(!D !C B A)+(!D C !B !A)+(!D C !B A)+(!D C B !A)+(!D C B A)), LSE_LINE_FILE_ID=3, LSE_LCOL=13, LSE_RCOL=44, LSE_LLINE=32, LSE_RLINE=32 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(11[2:53])
    defparam I1.init = 16'b0000000011111111;
    
endmodule
//
// Verilog Description of module inverter_U202
//

module inverter_U202 (\notGate[816]_keep , \notGate[817] ) /* synthesis syn_module_defined=1 */ ;
    input \notGate[816]_keep ;
    output \notGate[817] ;
    
    wire \notGate[816]_keep  /* synthesis alspreserve=1 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(25[15:22])
    
    LUT4 I1 (.A(\notGate[816]_keep ), .B(\notGate[816]_keep ), .C(\notGate[816]_keep ), 
         .D(\notGate[816]_keep ), .Z(\notGate[817] )) /* synthesis syn_instantiated=1, lut_function=((!D !C !B !A)+(!D !C !B A)+(!D !C B !A)+(!D !C B A)+(!D C !B !A)+(!D C !B A)+(!D C B !A)+(!D C B A)), LSE_LINE_FILE_ID=3, LSE_LCOL=13, LSE_RCOL=44, LSE_LLINE=32, LSE_RLINE=32 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(11[2:53])
    defparam I1.init = 16'b0000000011111111;
    
endmodule
//
// Verilog Description of module inverter_U203
//

module inverter_U203 (\notGate[815]_keep , \notGate[816] ) /* synthesis syn_module_defined=1 */ ;
    input \notGate[815]_keep ;
    output \notGate[816] ;
    
    wire \notGate[815]_keep  /* synthesis alspreserve=1 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(25[15:22])
    
    LUT4 I1 (.A(\notGate[815]_keep ), .B(\notGate[815]_keep ), .C(\notGate[815]_keep ), 
         .D(\notGate[815]_keep ), .Z(\notGate[816] )) /* synthesis syn_instantiated=1, lut_function=((!D !C !B !A)+(!D !C !B A)+(!D !C B !A)+(!D !C B A)+(!D C !B !A)+(!D C !B A)+(!D C B !A)+(!D C B A)), LSE_LINE_FILE_ID=3, LSE_LCOL=13, LSE_RCOL=44, LSE_LLINE=32, LSE_RLINE=32 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(11[2:53])
    defparam I1.init = 16'b0000000011111111;
    
endmodule
//
// Verilog Description of module inverter_U204
//

module inverter_U204 (\notGate[814]_keep , \notGate[815] ) /* synthesis syn_module_defined=1 */ ;
    input \notGate[814]_keep ;
    output \notGate[815] ;
    
    wire \notGate[814]_keep  /* synthesis alspreserve=1 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(25[15:22])
    
    LUT4 I1 (.A(\notGate[814]_keep ), .B(\notGate[814]_keep ), .C(\notGate[814]_keep ), 
         .D(\notGate[814]_keep ), .Z(\notGate[815] )) /* synthesis syn_instantiated=1, lut_function=((!D !C !B !A)+(!D !C !B A)+(!D !C B !A)+(!D !C B A)+(!D C !B !A)+(!D C !B A)+(!D C B !A)+(!D C B A)), LSE_LINE_FILE_ID=3, LSE_LCOL=13, LSE_RCOL=44, LSE_LLINE=32, LSE_RLINE=32 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(11[2:53])
    defparam I1.init = 16'b0000000011111111;
    
endmodule
//
// Verilog Description of module inverter_U205
//

module inverter_U205 (\notGate[813]_keep , \notGate[814] ) /* synthesis syn_module_defined=1 */ ;
    input \notGate[813]_keep ;
    output \notGate[814] ;
    
    wire \notGate[813]_keep  /* synthesis alspreserve=1 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(25[15:22])
    
    LUT4 I1 (.A(\notGate[813]_keep ), .B(\notGate[813]_keep ), .C(\notGate[813]_keep ), 
         .D(\notGate[813]_keep ), .Z(\notGate[814] )) /* synthesis syn_instantiated=1, lut_function=((!D !C !B !A)+(!D !C !B A)+(!D !C B !A)+(!D !C B A)+(!D C !B !A)+(!D C !B A)+(!D C B !A)+(!D C B A)), LSE_LINE_FILE_ID=3, LSE_LCOL=13, LSE_RCOL=44, LSE_LLINE=32, LSE_RLINE=32 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(11[2:53])
    defparam I1.init = 16'b0000000011111111;
    
endmodule
//
// Verilog Description of module inverter_U206
//

module inverter_U206 (\notGate[812]_keep , \notGate[813] ) /* synthesis syn_module_defined=1 */ ;
    input \notGate[812]_keep ;
    output \notGate[813] ;
    
    wire \notGate[812]_keep  /* synthesis alspreserve=1 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(25[15:22])
    
    LUT4 I1 (.A(\notGate[812]_keep ), .B(\notGate[812]_keep ), .C(\notGate[812]_keep ), 
         .D(\notGate[812]_keep ), .Z(\notGate[813] )) /* synthesis syn_instantiated=1, lut_function=((!D !C !B !A)+(!D !C !B A)+(!D !C B !A)+(!D !C B A)+(!D C !B !A)+(!D C !B A)+(!D C B !A)+(!D C B A)), LSE_LINE_FILE_ID=3, LSE_LCOL=13, LSE_RCOL=44, LSE_LLINE=32, LSE_RLINE=32 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(11[2:53])
    defparam I1.init = 16'b0000000011111111;
    
endmodule
//
// Verilog Description of module inverter_U207
//

module inverter_U207 (\notGate[811]_keep , \notGate[812] ) /* synthesis syn_module_defined=1 */ ;
    input \notGate[811]_keep ;
    output \notGate[812] ;
    
    wire \notGate[811]_keep  /* synthesis alspreserve=1 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(25[15:22])
    
    LUT4 I1 (.A(\notGate[811]_keep ), .B(\notGate[811]_keep ), .C(\notGate[811]_keep ), 
         .D(\notGate[811]_keep ), .Z(\notGate[812] )) /* synthesis syn_instantiated=1, lut_function=((!D !C !B !A)+(!D !C !B A)+(!D !C B !A)+(!D !C B A)+(!D C !B !A)+(!D C !B A)+(!D C B !A)+(!D C B A)), LSE_LINE_FILE_ID=3, LSE_LCOL=13, LSE_RCOL=44, LSE_LLINE=32, LSE_RLINE=32 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(11[2:53])
    defparam I1.init = 16'b0000000011111111;
    
endmodule
//
// Verilog Description of module inverter_U208
//

module inverter_U208 (\notGate[810]_keep , \notGate[811] ) /* synthesis syn_module_defined=1 */ ;
    input \notGate[810]_keep ;
    output \notGate[811] ;
    
    wire \notGate[810]_keep  /* synthesis alspreserve=1 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(25[15:22])
    
    LUT4 I1 (.A(\notGate[810]_keep ), .B(\notGate[810]_keep ), .C(\notGate[810]_keep ), 
         .D(\notGate[810]_keep ), .Z(\notGate[811] )) /* synthesis syn_instantiated=1, lut_function=((!D !C !B !A)+(!D !C !B A)+(!D !C B !A)+(!D !C B A)+(!D C !B !A)+(!D C !B A)+(!D C B !A)+(!D C B A)), LSE_LINE_FILE_ID=3, LSE_LCOL=13, LSE_RCOL=44, LSE_LLINE=32, LSE_RLINE=32 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(11[2:53])
    defparam I1.init = 16'b0000000011111111;
    
endmodule
//
// Verilog Description of module inverter_U209
//

module inverter_U209 (\notGate[809]_keep , \notGate[810] ) /* synthesis syn_module_defined=1 */ ;
    input \notGate[809]_keep ;
    output \notGate[810] ;
    
    wire \notGate[809]_keep  /* synthesis alspreserve=1 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(25[15:22])
    
    LUT4 I1 (.A(\notGate[809]_keep ), .B(\notGate[809]_keep ), .C(\notGate[809]_keep ), 
         .D(\notGate[809]_keep ), .Z(\notGate[810] )) /* synthesis syn_instantiated=1, lut_function=((!D !C !B !A)+(!D !C !B A)+(!D !C B !A)+(!D !C B A)+(!D C !B !A)+(!D C !B A)+(!D C B !A)+(!D C B A)), LSE_LINE_FILE_ID=3, LSE_LCOL=13, LSE_RCOL=44, LSE_LLINE=32, LSE_RLINE=32 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(11[2:53])
    defparam I1.init = 16'b0000000011111111;
    
endmodule
//
// Verilog Description of module inverter_U210
//

module inverter_U210 (\notGate[79]_keep , \notGate[80] ) /* synthesis syn_module_defined=1 */ ;
    input \notGate[79]_keep ;
    output \notGate[80] ;
    
    wire \notGate[79]_keep  /* synthesis alspreserve=1 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(25[15:22])
    
    LUT4 I1 (.A(\notGate[79]_keep ), .B(\notGate[79]_keep ), .C(\notGate[79]_keep ), 
         .D(\notGate[79]_keep ), .Z(\notGate[80] )) /* synthesis syn_instantiated=1, lut_function=((!D !C !B !A)+(!D !C !B A)+(!D !C B !A)+(!D !C B A)+(!D C !B !A)+(!D C !B A)+(!D C B !A)+(!D C B A)), LSE_LINE_FILE_ID=3, LSE_LCOL=13, LSE_RCOL=44, LSE_LLINE=32, LSE_RLINE=32 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(11[2:53])
    defparam I1.init = 16'b0000000011111111;
    
endmodule
//
// Verilog Description of module inverter_U211
//

module inverter_U211 (\notGate[808]_keep , \notGate[809] ) /* synthesis syn_module_defined=1 */ ;
    input \notGate[808]_keep ;
    output \notGate[809] ;
    
    wire \notGate[808]_keep  /* synthesis alspreserve=1 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(25[15:22])
    
    LUT4 I1 (.A(\notGate[808]_keep ), .B(\notGate[808]_keep ), .C(\notGate[808]_keep ), 
         .D(\notGate[808]_keep ), .Z(\notGate[809] )) /* synthesis syn_instantiated=1, lut_function=((!D !C !B !A)+(!D !C !B A)+(!D !C B !A)+(!D !C B A)+(!D C !B !A)+(!D C !B A)+(!D C B !A)+(!D C B A)), LSE_LINE_FILE_ID=3, LSE_LCOL=13, LSE_RCOL=44, LSE_LLINE=32, LSE_RLINE=32 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(11[2:53])
    defparam I1.init = 16'b0000000011111111;
    
endmodule
//
// Verilog Description of module inverter_U212
//

module inverter_U212 (\notGate[807]_keep , \notGate[808] ) /* synthesis syn_module_defined=1 */ ;
    input \notGate[807]_keep ;
    output \notGate[808] ;
    
    wire \notGate[807]_keep  /* synthesis alspreserve=1 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(25[15:22])
    
    LUT4 I1 (.A(\notGate[807]_keep ), .B(\notGate[807]_keep ), .C(\notGate[807]_keep ), 
         .D(\notGate[807]_keep ), .Z(\notGate[808] )) /* synthesis syn_instantiated=1, lut_function=((!D !C !B !A)+(!D !C !B A)+(!D !C B !A)+(!D !C B A)+(!D C !B !A)+(!D C !B A)+(!D C B !A)+(!D C B A)), LSE_LINE_FILE_ID=3, LSE_LCOL=13, LSE_RCOL=44, LSE_LLINE=32, LSE_RLINE=32 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(11[2:53])
    defparam I1.init = 16'b0000000011111111;
    
endmodule
//
// Verilog Description of module inverter_U213
//

module inverter_U213 (\notGate[806]_keep , \notGate[807] ) /* synthesis syn_module_defined=1 */ ;
    input \notGate[806]_keep ;
    output \notGate[807] ;
    
    wire \notGate[806]_keep  /* synthesis alspreserve=1 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(25[15:22])
    
    LUT4 I1 (.A(\notGate[806]_keep ), .B(\notGate[806]_keep ), .C(\notGate[806]_keep ), 
         .D(\notGate[806]_keep ), .Z(\notGate[807] )) /* synthesis syn_instantiated=1, lut_function=((!D !C !B !A)+(!D !C !B A)+(!D !C B !A)+(!D !C B A)+(!D C !B !A)+(!D C !B A)+(!D C B !A)+(!D C B A)), LSE_LINE_FILE_ID=3, LSE_LCOL=13, LSE_RCOL=44, LSE_LLINE=32, LSE_RLINE=32 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(11[2:53])
    defparam I1.init = 16'b0000000011111111;
    
endmodule
//
// Verilog Description of module inverter_U214
//

module inverter_U214 (\notGate[805]_keep , \notGate[806] ) /* synthesis syn_module_defined=1 */ ;
    input \notGate[805]_keep ;
    output \notGate[806] ;
    
    wire \notGate[805]_keep  /* synthesis alspreserve=1 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(25[15:22])
    
    LUT4 I1 (.A(\notGate[805]_keep ), .B(\notGate[805]_keep ), .C(\notGate[805]_keep ), 
         .D(\notGate[805]_keep ), .Z(\notGate[806] )) /* synthesis syn_instantiated=1, lut_function=((!D !C !B !A)+(!D !C !B A)+(!D !C B !A)+(!D !C B A)+(!D C !B !A)+(!D C !B A)+(!D C B !A)+(!D C B A)), LSE_LINE_FILE_ID=3, LSE_LCOL=13, LSE_RCOL=44, LSE_LLINE=32, LSE_RLINE=32 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(11[2:53])
    defparam I1.init = 16'b0000000011111111;
    
endmodule
//
// Verilog Description of module inverter_U215
//

module inverter_U215 (\notGate[804]_keep , \notGate[805] ) /* synthesis syn_module_defined=1 */ ;
    input \notGate[804]_keep ;
    output \notGate[805] ;
    
    wire \notGate[804]_keep  /* synthesis alspreserve=1 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(25[15:22])
    
    LUT4 I1 (.A(\notGate[804]_keep ), .B(\notGate[804]_keep ), .C(\notGate[804]_keep ), 
         .D(\notGate[804]_keep ), .Z(\notGate[805] )) /* synthesis syn_instantiated=1, lut_function=((!D !C !B !A)+(!D !C !B A)+(!D !C B !A)+(!D !C B A)+(!D C !B !A)+(!D C !B A)+(!D C B !A)+(!D C B A)), LSE_LINE_FILE_ID=3, LSE_LCOL=13, LSE_RCOL=44, LSE_LLINE=32, LSE_RLINE=32 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(11[2:53])
    defparam I1.init = 16'b0000000011111111;
    
endmodule
//
// Verilog Description of module inverter_U216
//

module inverter_U216 (\notGate[803]_keep , \notGate[804] ) /* synthesis syn_module_defined=1 */ ;
    input \notGate[803]_keep ;
    output \notGate[804] ;
    
    wire \notGate[803]_keep  /* synthesis alspreserve=1 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(25[15:22])
    
    LUT4 I1 (.A(\notGate[803]_keep ), .B(\notGate[803]_keep ), .C(\notGate[803]_keep ), 
         .D(\notGate[803]_keep ), .Z(\notGate[804] )) /* synthesis syn_instantiated=1, lut_function=((!D !C !B !A)+(!D !C !B A)+(!D !C B !A)+(!D !C B A)+(!D C !B !A)+(!D C !B A)+(!D C B !A)+(!D C B A)), LSE_LINE_FILE_ID=3, LSE_LCOL=13, LSE_RCOL=44, LSE_LLINE=32, LSE_RLINE=32 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(11[2:53])
    defparam I1.init = 16'b0000000011111111;
    
endmodule
//
// Verilog Description of module inverter_U217
//

module inverter_U217 (\notGate[802]_keep , \notGate[803] ) /* synthesis syn_module_defined=1 */ ;
    input \notGate[802]_keep ;
    output \notGate[803] ;
    
    wire \notGate[802]_keep  /* synthesis alspreserve=1 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(25[15:22])
    
    LUT4 I1 (.A(\notGate[802]_keep ), .B(\notGate[802]_keep ), .C(\notGate[802]_keep ), 
         .D(\notGate[802]_keep ), .Z(\notGate[803] )) /* synthesis syn_instantiated=1, lut_function=((!D !C !B !A)+(!D !C !B A)+(!D !C B !A)+(!D !C B A)+(!D C !B !A)+(!D C !B A)+(!D C B !A)+(!D C B A)), LSE_LINE_FILE_ID=3, LSE_LCOL=13, LSE_RCOL=44, LSE_LLINE=32, LSE_RLINE=32 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(11[2:53])
    defparam I1.init = 16'b0000000011111111;
    
endmodule
//
// Verilog Description of module inverter_U218
//

module inverter_U218 (\notGate[801]_keep , \notGate[802] ) /* synthesis syn_module_defined=1 */ ;
    input \notGate[801]_keep ;
    output \notGate[802] ;
    
    wire \notGate[801]_keep  /* synthesis alspreserve=1 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(25[15:22])
    
    LUT4 I1 (.A(\notGate[801]_keep ), .B(\notGate[801]_keep ), .C(\notGate[801]_keep ), 
         .D(\notGate[801]_keep ), .Z(\notGate[802] )) /* synthesis syn_instantiated=1, lut_function=((!D !C !B !A)+(!D !C !B A)+(!D !C B !A)+(!D !C B A)+(!D C !B !A)+(!D C !B A)+(!D C B !A)+(!D C B A)), LSE_LINE_FILE_ID=3, LSE_LCOL=13, LSE_RCOL=44, LSE_LLINE=32, LSE_RLINE=32 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(11[2:53])
    defparam I1.init = 16'b0000000011111111;
    
endmodule
//
// Verilog Description of module inverter_U219
//

module inverter_U219 (\notGate[800]_keep , \notGate[801] ) /* synthesis syn_module_defined=1 */ ;
    input \notGate[800]_keep ;
    output \notGate[801] ;
    
    wire \notGate[800]_keep  /* synthesis alspreserve=1 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(25[15:22])
    
    LUT4 I1 (.A(\notGate[800]_keep ), .B(\notGate[800]_keep ), .C(\notGate[800]_keep ), 
         .D(\notGate[800]_keep ), .Z(\notGate[801] )) /* synthesis syn_instantiated=1, lut_function=((!D !C !B !A)+(!D !C !B A)+(!D !C B !A)+(!D !C B A)+(!D C !B !A)+(!D C !B A)+(!D C B !A)+(!D C B A)), LSE_LINE_FILE_ID=3, LSE_LCOL=13, LSE_RCOL=44, LSE_LLINE=32, LSE_RLINE=32 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(11[2:53])
    defparam I1.init = 16'b0000000011111111;
    
endmodule
//
// Verilog Description of module inverter_U220
//

module inverter_U220 (\notGate[799]_keep , \notGate[800] ) /* synthesis syn_module_defined=1 */ ;
    input \notGate[799]_keep ;
    output \notGate[800] ;
    
    wire \notGate[799]_keep  /* synthesis alspreserve=1 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(25[15:22])
    
    LUT4 I1 (.A(\notGate[799]_keep ), .B(\notGate[799]_keep ), .C(\notGate[799]_keep ), 
         .D(\notGate[799]_keep ), .Z(\notGate[800] )) /* synthesis syn_instantiated=1, lut_function=((!D !C !B !A)+(!D !C !B A)+(!D !C B !A)+(!D !C B A)+(!D C !B !A)+(!D C !B A)+(!D C B !A)+(!D C B A)), LSE_LINE_FILE_ID=3, LSE_LCOL=13, LSE_RCOL=44, LSE_LLINE=32, LSE_RLINE=32 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(11[2:53])
    defparam I1.init = 16'b0000000011111111;
    
endmodule
//
// Verilog Description of module inverter_U221
//

module inverter_U221 (\notGate[6]_keep , \notGate[7] ) /* synthesis syn_module_defined=1 */ ;
    input \notGate[6]_keep ;
    output \notGate[7] ;
    
    wire \notGate[6]_keep  /* synthesis alspreserve=1 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(25[15:22])
    
    LUT4 I1 (.A(\notGate[6]_keep ), .B(\notGate[6]_keep ), .C(\notGate[6]_keep ), 
         .D(\notGate[6]_keep ), .Z(\notGate[7] )) /* synthesis syn_instantiated=1, lut_function=((!D !C !B !A)+(!D !C !B A)+(!D !C B !A)+(!D !C B A)+(!D C !B !A)+(!D C !B A)+(!D C B !A)+(!D C B A)), LSE_LINE_FILE_ID=3, LSE_LCOL=13, LSE_RCOL=44, LSE_LLINE=32, LSE_RLINE=32 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(11[2:53])
    defparam I1.init = 16'b0000000011111111;
    
endmodule
//
// Verilog Description of module inverter_U222
//

module inverter_U222 (\notGate[78]_keep , \notGate[79] ) /* synthesis syn_module_defined=1 */ ;
    input \notGate[78]_keep ;
    output \notGate[79] ;
    
    wire \notGate[78]_keep  /* synthesis alspreserve=1 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(25[15:22])
    
    LUT4 I1 (.A(\notGate[78]_keep ), .B(\notGate[78]_keep ), .C(\notGate[78]_keep ), 
         .D(\notGate[78]_keep ), .Z(\notGate[79] )) /* synthesis syn_instantiated=1, lut_function=((!D !C !B !A)+(!D !C !B A)+(!D !C B !A)+(!D !C B A)+(!D C !B !A)+(!D C !B A)+(!D C B !A)+(!D C B A)), LSE_LINE_FILE_ID=3, LSE_LCOL=13, LSE_RCOL=44, LSE_LLINE=32, LSE_RLINE=32 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(11[2:53])
    defparam I1.init = 16'b0000000011111111;
    
endmodule
//
// Verilog Description of module inverter_U223
//

module inverter_U223 (\notGate[798]_keep , \notGate[799] ) /* synthesis syn_module_defined=1 */ ;
    input \notGate[798]_keep ;
    output \notGate[799] ;
    
    wire \notGate[798]_keep  /* synthesis alspreserve=1 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(25[15:22])
    
    LUT4 I1 (.A(\notGate[798]_keep ), .B(\notGate[798]_keep ), .C(\notGate[798]_keep ), 
         .D(\notGate[798]_keep ), .Z(\notGate[799] )) /* synthesis syn_instantiated=1, lut_function=((!D !C !B !A)+(!D !C !B A)+(!D !C B !A)+(!D !C B A)+(!D C !B !A)+(!D C !B A)+(!D C B !A)+(!D C B A)), LSE_LINE_FILE_ID=3, LSE_LCOL=13, LSE_RCOL=44, LSE_LLINE=32, LSE_RLINE=32 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(11[2:53])
    defparam I1.init = 16'b0000000011111111;
    
endmodule
//
// Verilog Description of module inverter_U224
//

module inverter_U224 (\notGate[797]_keep , \notGate[798] ) /* synthesis syn_module_defined=1 */ ;
    input \notGate[797]_keep ;
    output \notGate[798] ;
    
    wire \notGate[797]_keep  /* synthesis alspreserve=1 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(25[15:22])
    
    LUT4 I1 (.A(\notGate[797]_keep ), .B(\notGate[797]_keep ), .C(\notGate[797]_keep ), 
         .D(\notGate[797]_keep ), .Z(\notGate[798] )) /* synthesis syn_instantiated=1, lut_function=((!D !C !B !A)+(!D !C !B A)+(!D !C B !A)+(!D !C B A)+(!D C !B !A)+(!D C !B A)+(!D C B !A)+(!D C B A)), LSE_LINE_FILE_ID=3, LSE_LCOL=13, LSE_RCOL=44, LSE_LLINE=32, LSE_RLINE=32 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(11[2:53])
    defparam I1.init = 16'b0000000011111111;
    
endmodule
//
// Verilog Description of module inverter_U225
//

module inverter_U225 (\notGate[796]_keep , \notGate[797] ) /* synthesis syn_module_defined=1 */ ;
    input \notGate[796]_keep ;
    output \notGate[797] ;
    
    wire \notGate[796]_keep  /* synthesis alspreserve=1 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(25[15:22])
    
    LUT4 I1 (.A(\notGate[796]_keep ), .B(\notGate[796]_keep ), .C(\notGate[796]_keep ), 
         .D(\notGate[796]_keep ), .Z(\notGate[797] )) /* synthesis syn_instantiated=1, lut_function=((!D !C !B !A)+(!D !C !B A)+(!D !C B !A)+(!D !C B A)+(!D C !B !A)+(!D C !B A)+(!D C B !A)+(!D C B A)), LSE_LINE_FILE_ID=3, LSE_LCOL=13, LSE_RCOL=44, LSE_LLINE=32, LSE_RLINE=32 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(11[2:53])
    defparam I1.init = 16'b0000000011111111;
    
endmodule
//
// Verilog Description of module inverter_U226
//

module inverter_U226 (\notGate[795]_keep , \notGate[796] ) /* synthesis syn_module_defined=1 */ ;
    input \notGate[795]_keep ;
    output \notGate[796] ;
    
    wire \notGate[795]_keep  /* synthesis alspreserve=1 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(25[15:22])
    
    LUT4 I1 (.A(\notGate[795]_keep ), .B(\notGate[795]_keep ), .C(\notGate[795]_keep ), 
         .D(\notGate[795]_keep ), .Z(\notGate[796] )) /* synthesis syn_instantiated=1, lut_function=((!D !C !B !A)+(!D !C !B A)+(!D !C B !A)+(!D !C B A)+(!D C !B !A)+(!D C !B A)+(!D C B !A)+(!D C B A)), LSE_LINE_FILE_ID=3, LSE_LCOL=13, LSE_RCOL=44, LSE_LLINE=32, LSE_RLINE=32 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(11[2:53])
    defparam I1.init = 16'b0000000011111111;
    
endmodule
//
// Verilog Description of module inverter_U227
//

module inverter_U227 (\notGate[794]_keep , \notGate[795] ) /* synthesis syn_module_defined=1 */ ;
    input \notGate[794]_keep ;
    output \notGate[795] ;
    
    wire \notGate[794]_keep  /* synthesis alspreserve=1 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(25[15:22])
    
    LUT4 I1 (.A(\notGate[794]_keep ), .B(\notGate[794]_keep ), .C(\notGate[794]_keep ), 
         .D(\notGate[794]_keep ), .Z(\notGate[795] )) /* synthesis syn_instantiated=1, lut_function=((!D !C !B !A)+(!D !C !B A)+(!D !C B !A)+(!D !C B A)+(!D C !B !A)+(!D C !B A)+(!D C B !A)+(!D C B A)), LSE_LINE_FILE_ID=3, LSE_LCOL=13, LSE_RCOL=44, LSE_LLINE=32, LSE_RLINE=32 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(11[2:53])
    defparam I1.init = 16'b0000000011111111;
    
endmodule
//
// Verilog Description of module inverter_U228
//

module inverter_U228 (\notGate[793]_keep , \notGate[794] ) /* synthesis syn_module_defined=1 */ ;
    input \notGate[793]_keep ;
    output \notGate[794] ;
    
    wire \notGate[793]_keep  /* synthesis alspreserve=1 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(25[15:22])
    
    LUT4 I1 (.A(\notGate[793]_keep ), .B(\notGate[793]_keep ), .C(\notGate[793]_keep ), 
         .D(\notGate[793]_keep ), .Z(\notGate[794] )) /* synthesis syn_instantiated=1, lut_function=((!D !C !B !A)+(!D !C !B A)+(!D !C B !A)+(!D !C B A)+(!D C !B !A)+(!D C !B A)+(!D C B !A)+(!D C B A)), LSE_LINE_FILE_ID=3, LSE_LCOL=13, LSE_RCOL=44, LSE_LLINE=32, LSE_RLINE=32 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(11[2:53])
    defparam I1.init = 16'b0000000011111111;
    
endmodule
//
// Verilog Description of module inverter_U229
//

module inverter_U229 (\notGate[792]_keep , \notGate[793] ) /* synthesis syn_module_defined=1 */ ;
    input \notGate[792]_keep ;
    output \notGate[793] ;
    
    wire \notGate[792]_keep  /* synthesis alspreserve=1 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(25[15:22])
    
    LUT4 I1 (.A(\notGate[792]_keep ), .B(\notGate[792]_keep ), .C(\notGate[792]_keep ), 
         .D(\notGate[792]_keep ), .Z(\notGate[793] )) /* synthesis syn_instantiated=1, lut_function=((!D !C !B !A)+(!D !C !B A)+(!D !C B !A)+(!D !C B A)+(!D C !B !A)+(!D C !B A)+(!D C B !A)+(!D C B A)), LSE_LINE_FILE_ID=3, LSE_LCOL=13, LSE_RCOL=44, LSE_LLINE=32, LSE_RLINE=32 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(11[2:53])
    defparam I1.init = 16'b0000000011111111;
    
endmodule
//
// Verilog Description of module inverter_U230
//

module inverter_U230 (\notGate[791]_keep , \notGate[792] ) /* synthesis syn_module_defined=1 */ ;
    input \notGate[791]_keep ;
    output \notGate[792] ;
    
    wire \notGate[791]_keep  /* synthesis alspreserve=1 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(25[15:22])
    
    LUT4 I1 (.A(\notGate[791]_keep ), .B(\notGate[791]_keep ), .C(\notGate[791]_keep ), 
         .D(\notGate[791]_keep ), .Z(\notGate[792] )) /* synthesis syn_instantiated=1, lut_function=((!D !C !B !A)+(!D !C !B A)+(!D !C B !A)+(!D !C B A)+(!D C !B !A)+(!D C !B A)+(!D C B !A)+(!D C B A)), LSE_LINE_FILE_ID=3, LSE_LCOL=13, LSE_RCOL=44, LSE_LLINE=32, LSE_RLINE=32 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(11[2:53])
    defparam I1.init = 16'b0000000011111111;
    
endmodule
//
// Verilog Description of module inverter_U231
//

module inverter_U231 (\notGate[790]_keep , \notGate[791] ) /* synthesis syn_module_defined=1 */ ;
    input \notGate[790]_keep ;
    output \notGate[791] ;
    
    wire \notGate[790]_keep  /* synthesis alspreserve=1 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(25[15:22])
    
    LUT4 I1 (.A(\notGate[790]_keep ), .B(\notGate[790]_keep ), .C(\notGate[790]_keep ), 
         .D(\notGate[790]_keep ), .Z(\notGate[791] )) /* synthesis syn_instantiated=1, lut_function=((!D !C !B !A)+(!D !C !B A)+(!D !C B !A)+(!D !C B A)+(!D C !B !A)+(!D C !B A)+(!D C B !A)+(!D C B A)), LSE_LINE_FILE_ID=3, LSE_LCOL=13, LSE_RCOL=44, LSE_LLINE=32, LSE_RLINE=32 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(11[2:53])
    defparam I1.init = 16'b0000000011111111;
    
endmodule
//
// Verilog Description of module inverter_U232
//

module inverter_U232 (\notGate[789]_keep , \notGate[790] ) /* synthesis syn_module_defined=1 */ ;
    input \notGate[789]_keep ;
    output \notGate[790] ;
    
    wire \notGate[789]_keep  /* synthesis alspreserve=1 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(25[15:22])
    
    LUT4 I1 (.A(\notGate[789]_keep ), .B(\notGate[789]_keep ), .C(\notGate[789]_keep ), 
         .D(\notGate[789]_keep ), .Z(\notGate[790] )) /* synthesis syn_instantiated=1, lut_function=((!D !C !B !A)+(!D !C !B A)+(!D !C B !A)+(!D !C B A)+(!D C !B !A)+(!D C !B A)+(!D C B !A)+(!D C B A)), LSE_LINE_FILE_ID=3, LSE_LCOL=13, LSE_RCOL=44, LSE_LLINE=32, LSE_RLINE=32 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(11[2:53])
    defparam I1.init = 16'b0000000011111111;
    
endmodule
//
// Verilog Description of module inverter_U233
//

module inverter_U233 (\notGate[77]_keep , \notGate[78] ) /* synthesis syn_module_defined=1 */ ;
    input \notGate[77]_keep ;
    output \notGate[78] ;
    
    wire \notGate[77]_keep  /* synthesis alspreserve=1 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(25[15:22])
    
    LUT4 I1 (.A(\notGate[77]_keep ), .B(\notGate[77]_keep ), .C(\notGate[77]_keep ), 
         .D(\notGate[77]_keep ), .Z(\notGate[78] )) /* synthesis syn_instantiated=1, lut_function=((!D !C !B !A)+(!D !C !B A)+(!D !C B !A)+(!D !C B A)+(!D C !B !A)+(!D C !B A)+(!D C B !A)+(!D C B A)), LSE_LINE_FILE_ID=3, LSE_LCOL=13, LSE_RCOL=44, LSE_LLINE=32, LSE_RLINE=32 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(11[2:53])
    defparam I1.init = 16'b0000000011111111;
    
endmodule
//
// Verilog Description of module inverter_U234
//

module inverter_U234 (\notGate[788]_keep , \notGate[789] ) /* synthesis syn_module_defined=1 */ ;
    input \notGate[788]_keep ;
    output \notGate[789] ;
    
    wire \notGate[788]_keep  /* synthesis alspreserve=1 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(25[15:22])
    
    LUT4 I1 (.A(\notGate[788]_keep ), .B(\notGate[788]_keep ), .C(\notGate[788]_keep ), 
         .D(\notGate[788]_keep ), .Z(\notGate[789] )) /* synthesis syn_instantiated=1, lut_function=((!D !C !B !A)+(!D !C !B A)+(!D !C B !A)+(!D !C B A)+(!D C !B !A)+(!D C !B A)+(!D C B !A)+(!D C B A)), LSE_LINE_FILE_ID=3, LSE_LCOL=13, LSE_RCOL=44, LSE_LLINE=32, LSE_RLINE=32 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(11[2:53])
    defparam I1.init = 16'b0000000011111111;
    
endmodule
//
// Verilog Description of module inverter_U235
//

module inverter_U235 (\notGate[787]_keep , \notGate[788] ) /* synthesis syn_module_defined=1 */ ;
    input \notGate[787]_keep ;
    output \notGate[788] ;
    
    wire \notGate[787]_keep  /* synthesis alspreserve=1 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(25[15:22])
    
    LUT4 I1 (.A(\notGate[787]_keep ), .B(\notGate[787]_keep ), .C(\notGate[787]_keep ), 
         .D(\notGate[787]_keep ), .Z(\notGate[788] )) /* synthesis syn_instantiated=1, lut_function=((!D !C !B !A)+(!D !C !B A)+(!D !C B !A)+(!D !C B A)+(!D C !B !A)+(!D C !B A)+(!D C B !A)+(!D C B A)), LSE_LINE_FILE_ID=3, LSE_LCOL=13, LSE_RCOL=44, LSE_LLINE=32, LSE_RLINE=32 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(11[2:53])
    defparam I1.init = 16'b0000000011111111;
    
endmodule
//
// Verilog Description of module inverter_U236
//

module inverter_U236 (\notGate[786]_keep , \notGate[787] ) /* synthesis syn_module_defined=1 */ ;
    input \notGate[786]_keep ;
    output \notGate[787] ;
    
    wire \notGate[786]_keep  /* synthesis alspreserve=1 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(25[15:22])
    
    LUT4 I1 (.A(\notGate[786]_keep ), .B(\notGate[786]_keep ), .C(\notGate[786]_keep ), 
         .D(\notGate[786]_keep ), .Z(\notGate[787] )) /* synthesis syn_instantiated=1, lut_function=((!D !C !B !A)+(!D !C !B A)+(!D !C B !A)+(!D !C B A)+(!D C !B !A)+(!D C !B A)+(!D C B !A)+(!D C B A)), LSE_LINE_FILE_ID=3, LSE_LCOL=13, LSE_RCOL=44, LSE_LLINE=32, LSE_RLINE=32 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(11[2:53])
    defparam I1.init = 16'b0000000011111111;
    
endmodule
//
// Verilog Description of module inverter_U237
//

module inverter_U237 (\notGate[785]_keep , \notGate[786] ) /* synthesis syn_module_defined=1 */ ;
    input \notGate[785]_keep ;
    output \notGate[786] ;
    
    wire \notGate[785]_keep  /* synthesis alspreserve=1 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(25[15:22])
    
    LUT4 I1 (.A(\notGate[785]_keep ), .B(\notGate[785]_keep ), .C(\notGate[785]_keep ), 
         .D(\notGate[785]_keep ), .Z(\notGate[786] )) /* synthesis syn_instantiated=1, lut_function=((!D !C !B !A)+(!D !C !B A)+(!D !C B !A)+(!D !C B A)+(!D C !B !A)+(!D C !B A)+(!D C B !A)+(!D C B A)), LSE_LINE_FILE_ID=3, LSE_LCOL=13, LSE_RCOL=44, LSE_LLINE=32, LSE_RLINE=32 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(11[2:53])
    defparam I1.init = 16'b0000000011111111;
    
endmodule
//
// Verilog Description of module inverter_U238
//

module inverter_U238 (\notGate[784]_keep , \notGate[785] ) /* synthesis syn_module_defined=1 */ ;
    input \notGate[784]_keep ;
    output \notGate[785] ;
    
    wire \notGate[784]_keep  /* synthesis alspreserve=1 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(25[15:22])
    
    LUT4 I1 (.A(\notGate[784]_keep ), .B(\notGate[784]_keep ), .C(\notGate[784]_keep ), 
         .D(\notGate[784]_keep ), .Z(\notGate[785] )) /* synthesis syn_instantiated=1, lut_function=((!D !C !B !A)+(!D !C !B A)+(!D !C B !A)+(!D !C B A)+(!D C !B !A)+(!D C !B A)+(!D C B !A)+(!D C B A)), LSE_LINE_FILE_ID=3, LSE_LCOL=13, LSE_RCOL=44, LSE_LLINE=32, LSE_RLINE=32 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(11[2:53])
    defparam I1.init = 16'b0000000011111111;
    
endmodule
//
// Verilog Description of module inverter_U239
//

module inverter_U239 (\notGate[783]_keep , \notGate[784] ) /* synthesis syn_module_defined=1 */ ;
    input \notGate[783]_keep ;
    output \notGate[784] ;
    
    wire \notGate[783]_keep  /* synthesis alspreserve=1 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(25[15:22])
    
    LUT4 I1 (.A(\notGate[783]_keep ), .B(\notGate[783]_keep ), .C(\notGate[783]_keep ), 
         .D(\notGate[783]_keep ), .Z(\notGate[784] )) /* synthesis syn_instantiated=1, lut_function=((!D !C !B !A)+(!D !C !B A)+(!D !C B !A)+(!D !C B A)+(!D C !B !A)+(!D C !B A)+(!D C B !A)+(!D C B A)), LSE_LINE_FILE_ID=3, LSE_LCOL=13, LSE_RCOL=44, LSE_LLINE=32, LSE_RLINE=32 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(11[2:53])
    defparam I1.init = 16'b0000000011111111;
    
endmodule
//
// Verilog Description of module inverter_U240
//

module inverter_U240 (\notGate[782]_keep , \notGate[783] ) /* synthesis syn_module_defined=1 */ ;
    input \notGate[782]_keep ;
    output \notGate[783] ;
    
    wire \notGate[782]_keep  /* synthesis alspreserve=1 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(25[15:22])
    
    LUT4 I1 (.A(\notGate[782]_keep ), .B(\notGate[782]_keep ), .C(\notGate[782]_keep ), 
         .D(\notGate[782]_keep ), .Z(\notGate[783] )) /* synthesis syn_instantiated=1, lut_function=((!D !C !B !A)+(!D !C !B A)+(!D !C B !A)+(!D !C B A)+(!D C !B !A)+(!D C !B A)+(!D C B !A)+(!D C B A)), LSE_LINE_FILE_ID=3, LSE_LCOL=13, LSE_RCOL=44, LSE_LLINE=32, LSE_RLINE=32 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(11[2:53])
    defparam I1.init = 16'b0000000011111111;
    
endmodule
//
// Verilog Description of module inverter_U241
//

module inverter_U241 (\notGate[781]_keep , \notGate[782] ) /* synthesis syn_module_defined=1 */ ;
    input \notGate[781]_keep ;
    output \notGate[782] ;
    
    wire \notGate[781]_keep  /* synthesis alspreserve=1 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(25[15:22])
    
    LUT4 I1 (.A(\notGate[781]_keep ), .B(\notGate[781]_keep ), .C(\notGate[781]_keep ), 
         .D(\notGate[781]_keep ), .Z(\notGate[782] )) /* synthesis syn_instantiated=1, lut_function=((!D !C !B !A)+(!D !C !B A)+(!D !C B !A)+(!D !C B A)+(!D C !B !A)+(!D C !B A)+(!D C B !A)+(!D C B A)), LSE_LINE_FILE_ID=3, LSE_LCOL=13, LSE_RCOL=44, LSE_LLINE=32, LSE_RLINE=32 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(11[2:53])
    defparam I1.init = 16'b0000000011111111;
    
endmodule
//
// Verilog Description of module inverter_U242
//

module inverter_U242 (\notGate[780]_keep , \notGate[781] ) /* synthesis syn_module_defined=1 */ ;
    input \notGate[780]_keep ;
    output \notGate[781] ;
    
    wire \notGate[780]_keep  /* synthesis alspreserve=1 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(25[15:22])
    
    LUT4 I1 (.A(\notGate[780]_keep ), .B(\notGate[780]_keep ), .C(\notGate[780]_keep ), 
         .D(\notGate[780]_keep ), .Z(\notGate[781] )) /* synthesis syn_instantiated=1, lut_function=((!D !C !B !A)+(!D !C !B A)+(!D !C B !A)+(!D !C B A)+(!D C !B !A)+(!D C !B A)+(!D C B !A)+(!D C B A)), LSE_LINE_FILE_ID=3, LSE_LCOL=13, LSE_RCOL=44, LSE_LLINE=32, LSE_RLINE=32 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(11[2:53])
    defparam I1.init = 16'b0000000011111111;
    
endmodule
//
// Verilog Description of module inverter_U243
//

module inverter_U243 (\notGate[779]_keep , \notGate[780] ) /* synthesis syn_module_defined=1 */ ;
    input \notGate[779]_keep ;
    output \notGate[780] ;
    
    wire \notGate[779]_keep  /* synthesis alspreserve=1 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(25[15:22])
    
    LUT4 I1 (.A(\notGate[779]_keep ), .B(\notGate[779]_keep ), .C(\notGate[779]_keep ), 
         .D(\notGate[779]_keep ), .Z(\notGate[780] )) /* synthesis syn_instantiated=1, lut_function=((!D !C !B !A)+(!D !C !B A)+(!D !C B !A)+(!D !C B A)+(!D C !B !A)+(!D C !B A)+(!D C B !A)+(!D C B A)), LSE_LINE_FILE_ID=3, LSE_LCOL=13, LSE_RCOL=44, LSE_LLINE=32, LSE_RLINE=32 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(11[2:53])
    defparam I1.init = 16'b0000000011111111;
    
endmodule
//
// Verilog Description of module inverter_U244
//

module inverter_U244 (\notGate[76]_keep , \notGate[77] ) /* synthesis syn_module_defined=1 */ ;
    input \notGate[76]_keep ;
    output \notGate[77] ;
    
    wire \notGate[76]_keep  /* synthesis alspreserve=1 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(25[15:22])
    
    LUT4 I1 (.A(\notGate[76]_keep ), .B(\notGate[76]_keep ), .C(\notGate[76]_keep ), 
         .D(\notGate[76]_keep ), .Z(\notGate[77] )) /* synthesis syn_instantiated=1, lut_function=((!D !C !B !A)+(!D !C !B A)+(!D !C B !A)+(!D !C B A)+(!D C !B !A)+(!D C !B A)+(!D C B !A)+(!D C B A)), LSE_LINE_FILE_ID=3, LSE_LCOL=13, LSE_RCOL=44, LSE_LLINE=32, LSE_RLINE=32 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(11[2:53])
    defparam I1.init = 16'b0000000011111111;
    
endmodule
//
// Verilog Description of module inverter_U245
//

module inverter_U245 (\notGate[778]_keep , \notGate[779] ) /* synthesis syn_module_defined=1 */ ;
    input \notGate[778]_keep ;
    output \notGate[779] ;
    
    wire \notGate[778]_keep  /* synthesis alspreserve=1 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(25[15:22])
    
    LUT4 I1 (.A(\notGate[778]_keep ), .B(\notGate[778]_keep ), .C(\notGate[778]_keep ), 
         .D(\notGate[778]_keep ), .Z(\notGate[779] )) /* synthesis syn_instantiated=1, lut_function=((!D !C !B !A)+(!D !C !B A)+(!D !C B !A)+(!D !C B A)+(!D C !B !A)+(!D C !B A)+(!D C B !A)+(!D C B A)), LSE_LINE_FILE_ID=3, LSE_LCOL=13, LSE_RCOL=44, LSE_LLINE=32, LSE_RLINE=32 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(11[2:53])
    defparam I1.init = 16'b0000000011111111;
    
endmodule
//
// Verilog Description of module inverter_U246
//

module inverter_U246 (\notGate[777]_keep , \notGate[778] ) /* synthesis syn_module_defined=1 */ ;
    input \notGate[777]_keep ;
    output \notGate[778] ;
    
    wire \notGate[777]_keep  /* synthesis alspreserve=1 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(25[15:22])
    
    LUT4 I1 (.A(\notGate[777]_keep ), .B(\notGate[777]_keep ), .C(\notGate[777]_keep ), 
         .D(\notGate[777]_keep ), .Z(\notGate[778] )) /* synthesis syn_instantiated=1, lut_function=((!D !C !B !A)+(!D !C !B A)+(!D !C B !A)+(!D !C B A)+(!D C !B !A)+(!D C !B A)+(!D C B !A)+(!D C B A)), LSE_LINE_FILE_ID=3, LSE_LCOL=13, LSE_RCOL=44, LSE_LLINE=32, LSE_RLINE=32 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(11[2:53])
    defparam I1.init = 16'b0000000011111111;
    
endmodule
//
// Verilog Description of module inverter_U247
//

module inverter_U247 (\notGate[776]_keep , \notGate[777] ) /* synthesis syn_module_defined=1 */ ;
    input \notGate[776]_keep ;
    output \notGate[777] ;
    
    wire \notGate[776]_keep  /* synthesis alspreserve=1 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(25[15:22])
    
    LUT4 I1 (.A(\notGate[776]_keep ), .B(\notGate[776]_keep ), .C(\notGate[776]_keep ), 
         .D(\notGate[776]_keep ), .Z(\notGate[777] )) /* synthesis syn_instantiated=1, lut_function=((!D !C !B !A)+(!D !C !B A)+(!D !C B !A)+(!D !C B A)+(!D C !B !A)+(!D C !B A)+(!D C B !A)+(!D C B A)), LSE_LINE_FILE_ID=3, LSE_LCOL=13, LSE_RCOL=44, LSE_LLINE=32, LSE_RLINE=32 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(11[2:53])
    defparam I1.init = 16'b0000000011111111;
    
endmodule
//
// Verilog Description of module inverter_U248
//

module inverter_U248 (\notGate[775]_keep , \notGate[776] ) /* synthesis syn_module_defined=1 */ ;
    input \notGate[775]_keep ;
    output \notGate[776] ;
    
    wire \notGate[775]_keep  /* synthesis alspreserve=1 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(25[15:22])
    
    LUT4 I1 (.A(\notGate[775]_keep ), .B(\notGate[775]_keep ), .C(\notGate[775]_keep ), 
         .D(\notGate[775]_keep ), .Z(\notGate[776] )) /* synthesis syn_instantiated=1, lut_function=((!D !C !B !A)+(!D !C !B A)+(!D !C B !A)+(!D !C B A)+(!D C !B !A)+(!D C !B A)+(!D C B !A)+(!D C B A)), LSE_LINE_FILE_ID=3, LSE_LCOL=13, LSE_RCOL=44, LSE_LLINE=32, LSE_RLINE=32 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(11[2:53])
    defparam I1.init = 16'b0000000011111111;
    
endmodule
//
// Verilog Description of module inverter_U249
//

module inverter_U249 (\notGate[774]_keep , \notGate[775] ) /* synthesis syn_module_defined=1 */ ;
    input \notGate[774]_keep ;
    output \notGate[775] ;
    
    wire \notGate[774]_keep  /* synthesis alspreserve=1 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(25[15:22])
    
    LUT4 I1 (.A(\notGate[774]_keep ), .B(\notGate[774]_keep ), .C(\notGate[774]_keep ), 
         .D(\notGate[774]_keep ), .Z(\notGate[775] )) /* synthesis syn_instantiated=1, lut_function=((!D !C !B !A)+(!D !C !B A)+(!D !C B !A)+(!D !C B A)+(!D C !B !A)+(!D C !B A)+(!D C B !A)+(!D C B A)), LSE_LINE_FILE_ID=3, LSE_LCOL=13, LSE_RCOL=44, LSE_LLINE=32, LSE_RLINE=32 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(11[2:53])
    defparam I1.init = 16'b0000000011111111;
    
endmodule
//
// Verilog Description of module inverter_U250
//

module inverter_U250 (\notGate[773]_keep , \notGate[774] ) /* synthesis syn_module_defined=1 */ ;
    input \notGate[773]_keep ;
    output \notGate[774] ;
    
    wire \notGate[773]_keep  /* synthesis alspreserve=1 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(25[15:22])
    
    LUT4 I1 (.A(\notGate[773]_keep ), .B(\notGate[773]_keep ), .C(\notGate[773]_keep ), 
         .D(\notGate[773]_keep ), .Z(\notGate[774] )) /* synthesis syn_instantiated=1, lut_function=((!D !C !B !A)+(!D !C !B A)+(!D !C B !A)+(!D !C B A)+(!D C !B !A)+(!D C !B A)+(!D C B !A)+(!D C B A)), LSE_LINE_FILE_ID=3, LSE_LCOL=13, LSE_RCOL=44, LSE_LLINE=32, LSE_RLINE=32 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(11[2:53])
    defparam I1.init = 16'b0000000011111111;
    
endmodule
//
// Verilog Description of module inverter_U251
//

module inverter_U251 (\notGate[772]_keep , \notGate[773] ) /* synthesis syn_module_defined=1 */ ;
    input \notGate[772]_keep ;
    output \notGate[773] ;
    
    wire \notGate[772]_keep  /* synthesis alspreserve=1 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(25[15:22])
    
    LUT4 I1 (.A(\notGate[772]_keep ), .B(\notGate[772]_keep ), .C(\notGate[772]_keep ), 
         .D(\notGate[772]_keep ), .Z(\notGate[773] )) /* synthesis syn_instantiated=1, lut_function=((!D !C !B !A)+(!D !C !B A)+(!D !C B !A)+(!D !C B A)+(!D C !B !A)+(!D C !B A)+(!D C B !A)+(!D C B A)), LSE_LINE_FILE_ID=3, LSE_LCOL=13, LSE_RCOL=44, LSE_LLINE=32, LSE_RLINE=32 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(11[2:53])
    defparam I1.init = 16'b0000000011111111;
    
endmodule
//
// Verilog Description of module inverter_U252
//

module inverter_U252 (\notGate[771]_keep , \notGate[772] ) /* synthesis syn_module_defined=1 */ ;
    input \notGate[771]_keep ;
    output \notGate[772] ;
    
    wire \notGate[771]_keep  /* synthesis alspreserve=1 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(25[15:22])
    
    LUT4 I1 (.A(\notGate[771]_keep ), .B(\notGate[771]_keep ), .C(\notGate[771]_keep ), 
         .D(\notGate[771]_keep ), .Z(\notGate[772] )) /* synthesis syn_instantiated=1, lut_function=((!D !C !B !A)+(!D !C !B A)+(!D !C B !A)+(!D !C B A)+(!D C !B !A)+(!D C !B A)+(!D C B !A)+(!D C B A)), LSE_LINE_FILE_ID=3, LSE_LCOL=13, LSE_RCOL=44, LSE_LLINE=32, LSE_RLINE=32 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(11[2:53])
    defparam I1.init = 16'b0000000011111111;
    
endmodule
//
// Verilog Description of module inverter_U253
//

module inverter_U253 (\notGate[770]_keep , \notGate[771] ) /* synthesis syn_module_defined=1 */ ;
    input \notGate[770]_keep ;
    output \notGate[771] ;
    
    wire \notGate[770]_keep  /* synthesis alspreserve=1 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(25[15:22])
    
    LUT4 I1 (.A(\notGate[770]_keep ), .B(\notGate[770]_keep ), .C(\notGate[770]_keep ), 
         .D(\notGate[770]_keep ), .Z(\notGate[771] )) /* synthesis syn_instantiated=1, lut_function=((!D !C !B !A)+(!D !C !B A)+(!D !C B !A)+(!D !C B A)+(!D C !B !A)+(!D C !B A)+(!D C B !A)+(!D C B A)), LSE_LINE_FILE_ID=3, LSE_LCOL=13, LSE_RCOL=44, LSE_LLINE=32, LSE_RLINE=32 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(11[2:53])
    defparam I1.init = 16'b0000000011111111;
    
endmodule
//
// Verilog Description of module inverter_U254
//

module inverter_U254 (\notGate[769]_keep , \notGate[770] ) /* synthesis syn_module_defined=1 */ ;
    input \notGate[769]_keep ;
    output \notGate[770] ;
    
    wire \notGate[769]_keep  /* synthesis alspreserve=1 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(25[15:22])
    
    LUT4 I1 (.A(\notGate[769]_keep ), .B(\notGate[769]_keep ), .C(\notGate[769]_keep ), 
         .D(\notGate[769]_keep ), .Z(\notGate[770] )) /* synthesis syn_instantiated=1, lut_function=((!D !C !B !A)+(!D !C !B A)+(!D !C B !A)+(!D !C B A)+(!D C !B !A)+(!D C !B A)+(!D C B !A)+(!D C B A)), LSE_LINE_FILE_ID=3, LSE_LCOL=13, LSE_RCOL=44, LSE_LLINE=32, LSE_RLINE=32 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(11[2:53])
    defparam I1.init = 16'b0000000011111111;
    
endmodule
//
// Verilog Description of module inverter_U255
//

module inverter_U255 (\notGate[75]_keep , \notGate[76] ) /* synthesis syn_module_defined=1 */ ;
    input \notGate[75]_keep ;
    output \notGate[76] ;
    
    wire \notGate[75]_keep  /* synthesis alspreserve=1 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(25[15:22])
    
    LUT4 I1 (.A(\notGate[75]_keep ), .B(\notGate[75]_keep ), .C(\notGate[75]_keep ), 
         .D(\notGate[75]_keep ), .Z(\notGate[76] )) /* synthesis syn_instantiated=1, lut_function=((!D !C !B !A)+(!D !C !B A)+(!D !C B !A)+(!D !C B A)+(!D C !B !A)+(!D C !B A)+(!D C B !A)+(!D C B A)), LSE_LINE_FILE_ID=3, LSE_LCOL=13, LSE_RCOL=44, LSE_LLINE=32, LSE_RLINE=32 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(11[2:53])
    defparam I1.init = 16'b0000000011111111;
    
endmodule
//
// Verilog Description of module inverter_U256
//

module inverter_U256 (\notGate[768]_keep , \notGate[769] ) /* synthesis syn_module_defined=1 */ ;
    input \notGate[768]_keep ;
    output \notGate[769] ;
    
    wire \notGate[768]_keep  /* synthesis alspreserve=1 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(25[15:22])
    
    LUT4 I1 (.A(\notGate[768]_keep ), .B(\notGate[768]_keep ), .C(\notGate[768]_keep ), 
         .D(\notGate[768]_keep ), .Z(\notGate[769] )) /* synthesis syn_instantiated=1, lut_function=((!D !C !B !A)+(!D !C !B A)+(!D !C B !A)+(!D !C B A)+(!D C !B !A)+(!D C !B A)+(!D C B !A)+(!D C B A)), LSE_LINE_FILE_ID=3, LSE_LCOL=13, LSE_RCOL=44, LSE_LLINE=32, LSE_RLINE=32 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(11[2:53])
    defparam I1.init = 16'b0000000011111111;
    
endmodule
//
// Verilog Description of module inverter_U257
//

module inverter_U257 (\notGate[767]_keep , \notGate[768] ) /* synthesis syn_module_defined=1 */ ;
    input \notGate[767]_keep ;
    output \notGate[768] ;
    
    wire \notGate[767]_keep  /* synthesis alspreserve=1 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(25[15:22])
    
    LUT4 I1 (.A(\notGate[767]_keep ), .B(\notGate[767]_keep ), .C(\notGate[767]_keep ), 
         .D(\notGate[767]_keep ), .Z(\notGate[768] )) /* synthesis syn_instantiated=1, lut_function=((!D !C !B !A)+(!D !C !B A)+(!D !C B !A)+(!D !C B A)+(!D C !B !A)+(!D C !B A)+(!D C B !A)+(!D C B A)), LSE_LINE_FILE_ID=3, LSE_LCOL=13, LSE_RCOL=44, LSE_LLINE=32, LSE_RLINE=32 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(11[2:53])
    defparam I1.init = 16'b0000000011111111;
    
endmodule
//
// Verilog Description of module inverter_U258
//

module inverter_U258 (\notGate[766]_keep , \notGate[767] ) /* synthesis syn_module_defined=1 */ ;
    input \notGate[766]_keep ;
    output \notGate[767] ;
    
    wire \notGate[766]_keep  /* synthesis alspreserve=1 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(25[15:22])
    
    LUT4 I1 (.A(\notGate[766]_keep ), .B(\notGate[766]_keep ), .C(\notGate[766]_keep ), 
         .D(\notGate[766]_keep ), .Z(\notGate[767] )) /* synthesis syn_instantiated=1, lut_function=((!D !C !B !A)+(!D !C !B A)+(!D !C B !A)+(!D !C B A)+(!D C !B !A)+(!D C !B A)+(!D C B !A)+(!D C B A)), LSE_LINE_FILE_ID=3, LSE_LCOL=13, LSE_RCOL=44, LSE_LLINE=32, LSE_RLINE=32 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(11[2:53])
    defparam I1.init = 16'b0000000011111111;
    
endmodule
//
// Verilog Description of module inverter_U259
//

module inverter_U259 (\notGate[765]_keep , \notGate[766] ) /* synthesis syn_module_defined=1 */ ;
    input \notGate[765]_keep ;
    output \notGate[766] ;
    
    wire \notGate[765]_keep  /* synthesis alspreserve=1 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(25[15:22])
    
    LUT4 I1 (.A(\notGate[765]_keep ), .B(\notGate[765]_keep ), .C(\notGate[765]_keep ), 
         .D(\notGate[765]_keep ), .Z(\notGate[766] )) /* synthesis syn_instantiated=1, lut_function=((!D !C !B !A)+(!D !C !B A)+(!D !C B !A)+(!D !C B A)+(!D C !B !A)+(!D C !B A)+(!D C B !A)+(!D C B A)), LSE_LINE_FILE_ID=3, LSE_LCOL=13, LSE_RCOL=44, LSE_LLINE=32, LSE_RLINE=32 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(11[2:53])
    defparam I1.init = 16'b0000000011111111;
    
endmodule
//
// Verilog Description of module inverter_U260
//

module inverter_U260 (\notGate[764]_keep , \notGate[765] ) /* synthesis syn_module_defined=1 */ ;
    input \notGate[764]_keep ;
    output \notGate[765] ;
    
    wire \notGate[764]_keep  /* synthesis alspreserve=1 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(25[15:22])
    
    LUT4 I1 (.A(\notGate[764]_keep ), .B(\notGate[764]_keep ), .C(\notGate[764]_keep ), 
         .D(\notGate[764]_keep ), .Z(\notGate[765] )) /* synthesis syn_instantiated=1, lut_function=((!D !C !B !A)+(!D !C !B A)+(!D !C B !A)+(!D !C B A)+(!D C !B !A)+(!D C !B A)+(!D C B !A)+(!D C B A)), LSE_LINE_FILE_ID=3, LSE_LCOL=13, LSE_RCOL=44, LSE_LLINE=32, LSE_RLINE=32 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(11[2:53])
    defparam I1.init = 16'b0000000011111111;
    
endmodule
//
// Verilog Description of module inverter_U261
//

module inverter_U261 (\notGate[763]_keep , \notGate[764] ) /* synthesis syn_module_defined=1 */ ;
    input \notGate[763]_keep ;
    output \notGate[764] ;
    
    wire \notGate[763]_keep  /* synthesis alspreserve=1 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(25[15:22])
    
    LUT4 I1 (.A(\notGate[763]_keep ), .B(\notGate[763]_keep ), .C(\notGate[763]_keep ), 
         .D(\notGate[763]_keep ), .Z(\notGate[764] )) /* synthesis syn_instantiated=1, lut_function=((!D !C !B !A)+(!D !C !B A)+(!D !C B !A)+(!D !C B A)+(!D C !B !A)+(!D C !B A)+(!D C B !A)+(!D C B A)), LSE_LINE_FILE_ID=3, LSE_LCOL=13, LSE_RCOL=44, LSE_LLINE=32, LSE_RLINE=32 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(11[2:53])
    defparam I1.init = 16'b0000000011111111;
    
endmodule
//
// Verilog Description of module inverter_U262
//

module inverter_U262 (\notGate[762]_keep , \notGate[763] ) /* synthesis syn_module_defined=1 */ ;
    input \notGate[762]_keep ;
    output \notGate[763] ;
    
    wire \notGate[762]_keep  /* synthesis alspreserve=1 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(25[15:22])
    
    LUT4 I1 (.A(\notGate[762]_keep ), .B(\notGate[762]_keep ), .C(\notGate[762]_keep ), 
         .D(\notGate[762]_keep ), .Z(\notGate[763] )) /* synthesis syn_instantiated=1, lut_function=((!D !C !B !A)+(!D !C !B A)+(!D !C B !A)+(!D !C B A)+(!D C !B !A)+(!D C !B A)+(!D C B !A)+(!D C B A)), LSE_LINE_FILE_ID=3, LSE_LCOL=13, LSE_RCOL=44, LSE_LLINE=32, LSE_RLINE=32 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(11[2:53])
    defparam I1.init = 16'b0000000011111111;
    
endmodule
//
// Verilog Description of module inverter_U263
//

module inverter_U263 (\notGate[761]_keep , \notGate[762] ) /* synthesis syn_module_defined=1 */ ;
    input \notGate[761]_keep ;
    output \notGate[762] ;
    
    wire \notGate[761]_keep  /* synthesis alspreserve=1 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(25[15:22])
    
    LUT4 I1 (.A(\notGate[761]_keep ), .B(\notGate[761]_keep ), .C(\notGate[761]_keep ), 
         .D(\notGate[761]_keep ), .Z(\notGate[762] )) /* synthesis syn_instantiated=1, lut_function=((!D !C !B !A)+(!D !C !B A)+(!D !C B !A)+(!D !C B A)+(!D C !B !A)+(!D C !B A)+(!D C B !A)+(!D C B A)), LSE_LINE_FILE_ID=3, LSE_LCOL=13, LSE_RCOL=44, LSE_LLINE=32, LSE_RLINE=32 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(11[2:53])
    defparam I1.init = 16'b0000000011111111;
    
endmodule
//
// Verilog Description of module inverter_U264
//

module inverter_U264 (\notGate[760]_keep , \notGate[761] ) /* synthesis syn_module_defined=1 */ ;
    input \notGate[760]_keep ;
    output \notGate[761] ;
    
    wire \notGate[760]_keep  /* synthesis alspreserve=1 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(25[15:22])
    
    LUT4 I1 (.A(\notGate[760]_keep ), .B(\notGate[760]_keep ), .C(\notGate[760]_keep ), 
         .D(\notGate[760]_keep ), .Z(\notGate[761] )) /* synthesis syn_instantiated=1, lut_function=((!D !C !B !A)+(!D !C !B A)+(!D !C B !A)+(!D !C B A)+(!D C !B !A)+(!D C !B A)+(!D C B !A)+(!D C B A)), LSE_LINE_FILE_ID=3, LSE_LCOL=13, LSE_RCOL=44, LSE_LLINE=32, LSE_RLINE=32 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(11[2:53])
    defparam I1.init = 16'b0000000011111111;
    
endmodule
//
// Verilog Description of module inverter_U265
//

module inverter_U265 (\notGate[759]_keep , \notGate[760] ) /* synthesis syn_module_defined=1 */ ;
    input \notGate[759]_keep ;
    output \notGate[760] ;
    
    wire \notGate[759]_keep  /* synthesis alspreserve=1 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(25[15:22])
    
    LUT4 I1 (.A(\notGate[759]_keep ), .B(\notGate[759]_keep ), .C(\notGate[759]_keep ), 
         .D(\notGate[759]_keep ), .Z(\notGate[760] )) /* synthesis syn_instantiated=1, lut_function=((!D !C !B !A)+(!D !C !B A)+(!D !C B !A)+(!D !C B A)+(!D C !B !A)+(!D C !B A)+(!D C B !A)+(!D C B A)), LSE_LINE_FILE_ID=3, LSE_LCOL=13, LSE_RCOL=44, LSE_LLINE=32, LSE_RLINE=32 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(11[2:53])
    defparam I1.init = 16'b0000000011111111;
    
endmodule
//
// Verilog Description of module inverter_U266
//

module inverter_U266 (\notGate[74]_keep , \notGate[75] ) /* synthesis syn_module_defined=1 */ ;
    input \notGate[74]_keep ;
    output \notGate[75] ;
    
    wire \notGate[74]_keep  /* synthesis alspreserve=1 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(25[15:22])
    
    LUT4 I1 (.A(\notGate[74]_keep ), .B(\notGate[74]_keep ), .C(\notGate[74]_keep ), 
         .D(\notGate[74]_keep ), .Z(\notGate[75] )) /* synthesis syn_instantiated=1, lut_function=((!D !C !B !A)+(!D !C !B A)+(!D !C B !A)+(!D !C B A)+(!D C !B !A)+(!D C !B A)+(!D C B !A)+(!D C B A)), LSE_LINE_FILE_ID=3, LSE_LCOL=13, LSE_RCOL=44, LSE_LLINE=32, LSE_RLINE=32 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(11[2:53])
    defparam I1.init = 16'b0000000011111111;
    
endmodule
//
// Verilog Description of module inverter_U267
//

module inverter_U267 (\notGate[758]_keep , \notGate[759] ) /* synthesis syn_module_defined=1 */ ;
    input \notGate[758]_keep ;
    output \notGate[759] ;
    
    wire \notGate[758]_keep  /* synthesis alspreserve=1 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(25[15:22])
    
    LUT4 I1 (.A(\notGate[758]_keep ), .B(\notGate[758]_keep ), .C(\notGate[758]_keep ), 
         .D(\notGate[758]_keep ), .Z(\notGate[759] )) /* synthesis syn_instantiated=1, lut_function=((!D !C !B !A)+(!D !C !B A)+(!D !C B !A)+(!D !C B A)+(!D C !B !A)+(!D C !B A)+(!D C B !A)+(!D C B A)), LSE_LINE_FILE_ID=3, LSE_LCOL=13, LSE_RCOL=44, LSE_LLINE=32, LSE_RLINE=32 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(11[2:53])
    defparam I1.init = 16'b0000000011111111;
    
endmodule
//
// Verilog Description of module inverter_U268
//

module inverter_U268 (\notGate[757]_keep , \notGate[758] ) /* synthesis syn_module_defined=1 */ ;
    input \notGate[757]_keep ;
    output \notGate[758] ;
    
    wire \notGate[757]_keep  /* synthesis alspreserve=1 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(25[15:22])
    
    LUT4 I1 (.A(\notGate[757]_keep ), .B(\notGate[757]_keep ), .C(\notGate[757]_keep ), 
         .D(\notGate[757]_keep ), .Z(\notGate[758] )) /* synthesis syn_instantiated=1, lut_function=((!D !C !B !A)+(!D !C !B A)+(!D !C B !A)+(!D !C B A)+(!D C !B !A)+(!D C !B A)+(!D C B !A)+(!D C B A)), LSE_LINE_FILE_ID=3, LSE_LCOL=13, LSE_RCOL=44, LSE_LLINE=32, LSE_RLINE=32 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(11[2:53])
    defparam I1.init = 16'b0000000011111111;
    
endmodule
//
// Verilog Description of module inverter_U269
//

module inverter_U269 (\notGate[756]_keep , \notGate[757] ) /* synthesis syn_module_defined=1 */ ;
    input \notGate[756]_keep ;
    output \notGate[757] ;
    
    wire \notGate[756]_keep  /* synthesis alspreserve=1 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(25[15:22])
    
    LUT4 I1 (.A(\notGate[756]_keep ), .B(\notGate[756]_keep ), .C(\notGate[756]_keep ), 
         .D(\notGate[756]_keep ), .Z(\notGate[757] )) /* synthesis syn_instantiated=1, lut_function=((!D !C !B !A)+(!D !C !B A)+(!D !C B !A)+(!D !C B A)+(!D C !B !A)+(!D C !B A)+(!D C B !A)+(!D C B A)), LSE_LINE_FILE_ID=3, LSE_LCOL=13, LSE_RCOL=44, LSE_LLINE=32, LSE_RLINE=32 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(11[2:53])
    defparam I1.init = 16'b0000000011111111;
    
endmodule
//
// Verilog Description of module inverter_U270
//

module inverter_U270 (\notGate[755]_keep , \notGate[756] ) /* synthesis syn_module_defined=1 */ ;
    input \notGate[755]_keep ;
    output \notGate[756] ;
    
    wire \notGate[755]_keep  /* synthesis alspreserve=1 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(25[15:22])
    
    LUT4 I1 (.A(\notGate[755]_keep ), .B(\notGate[755]_keep ), .C(\notGate[755]_keep ), 
         .D(\notGate[755]_keep ), .Z(\notGate[756] )) /* synthesis syn_instantiated=1, lut_function=((!D !C !B !A)+(!D !C !B A)+(!D !C B !A)+(!D !C B A)+(!D C !B !A)+(!D C !B A)+(!D C B !A)+(!D C B A)), LSE_LINE_FILE_ID=3, LSE_LCOL=13, LSE_RCOL=44, LSE_LLINE=32, LSE_RLINE=32 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(11[2:53])
    defparam I1.init = 16'b0000000011111111;
    
endmodule
//
// Verilog Description of module inverter_U271
//

module inverter_U271 (\notGate[754]_keep , \notGate[755] ) /* synthesis syn_module_defined=1 */ ;
    input \notGate[754]_keep ;
    output \notGate[755] ;
    
    wire \notGate[754]_keep  /* synthesis alspreserve=1 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(25[15:22])
    
    LUT4 I1 (.A(\notGate[754]_keep ), .B(\notGate[754]_keep ), .C(\notGate[754]_keep ), 
         .D(\notGate[754]_keep ), .Z(\notGate[755] )) /* synthesis syn_instantiated=1, lut_function=((!D !C !B !A)+(!D !C !B A)+(!D !C B !A)+(!D !C B A)+(!D C !B !A)+(!D C !B A)+(!D C B !A)+(!D C B A)), LSE_LINE_FILE_ID=3, LSE_LCOL=13, LSE_RCOL=44, LSE_LLINE=32, LSE_RLINE=32 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(11[2:53])
    defparam I1.init = 16'b0000000011111111;
    
endmodule
//
// Verilog Description of module inverter_U272
//

module inverter_U272 (\notGate[753]_keep , \notGate[754] ) /* synthesis syn_module_defined=1 */ ;
    input \notGate[753]_keep ;
    output \notGate[754] ;
    
    wire \notGate[753]_keep  /* synthesis alspreserve=1 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(25[15:22])
    
    LUT4 I1 (.A(\notGate[753]_keep ), .B(\notGate[753]_keep ), .C(\notGate[753]_keep ), 
         .D(\notGate[753]_keep ), .Z(\notGate[754] )) /* synthesis syn_instantiated=1, lut_function=((!D !C !B !A)+(!D !C !B A)+(!D !C B !A)+(!D !C B A)+(!D C !B !A)+(!D C !B A)+(!D C B !A)+(!D C B A)), LSE_LINE_FILE_ID=3, LSE_LCOL=13, LSE_RCOL=44, LSE_LLINE=32, LSE_RLINE=32 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(11[2:53])
    defparam I1.init = 16'b0000000011111111;
    
endmodule
//
// Verilog Description of module inverter_U273
//

module inverter_U273 (\notGate[752]_keep , \notGate[753] ) /* synthesis syn_module_defined=1 */ ;
    input \notGate[752]_keep ;
    output \notGate[753] ;
    
    wire \notGate[752]_keep  /* synthesis alspreserve=1 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(25[15:22])
    
    LUT4 I1 (.A(\notGate[752]_keep ), .B(\notGate[752]_keep ), .C(\notGate[752]_keep ), 
         .D(\notGate[752]_keep ), .Z(\notGate[753] )) /* synthesis syn_instantiated=1, lut_function=((!D !C !B !A)+(!D !C !B A)+(!D !C B !A)+(!D !C B A)+(!D C !B !A)+(!D C !B A)+(!D C B !A)+(!D C B A)), LSE_LINE_FILE_ID=3, LSE_LCOL=13, LSE_RCOL=44, LSE_LLINE=32, LSE_RLINE=32 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(11[2:53])
    defparam I1.init = 16'b0000000011111111;
    
endmodule
//
// Verilog Description of module inverter_U274
//

module inverter_U274 (\notGate[751]_keep , \notGate[752] ) /* synthesis syn_module_defined=1 */ ;
    input \notGate[751]_keep ;
    output \notGate[752] ;
    
    wire \notGate[751]_keep  /* synthesis alspreserve=1 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(25[15:22])
    
    LUT4 I1 (.A(\notGate[751]_keep ), .B(\notGate[751]_keep ), .C(\notGate[751]_keep ), 
         .D(\notGate[751]_keep ), .Z(\notGate[752] )) /* synthesis syn_instantiated=1, lut_function=((!D !C !B !A)+(!D !C !B A)+(!D !C B !A)+(!D !C B A)+(!D C !B !A)+(!D C !B A)+(!D C B !A)+(!D C B A)), LSE_LINE_FILE_ID=3, LSE_LCOL=13, LSE_RCOL=44, LSE_LLINE=32, LSE_RLINE=32 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(11[2:53])
    defparam I1.init = 16'b0000000011111111;
    
endmodule
//
// Verilog Description of module inverter_U275
//

module inverter_U275 (\notGate[750]_keep , \notGate[751] ) /* synthesis syn_module_defined=1 */ ;
    input \notGate[750]_keep ;
    output \notGate[751] ;
    
    wire \notGate[750]_keep  /* synthesis alspreserve=1 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(25[15:22])
    
    LUT4 I1 (.A(\notGate[750]_keep ), .B(\notGate[750]_keep ), .C(\notGate[750]_keep ), 
         .D(\notGate[750]_keep ), .Z(\notGate[751] )) /* synthesis syn_instantiated=1, lut_function=((!D !C !B !A)+(!D !C !B A)+(!D !C B !A)+(!D !C B A)+(!D C !B !A)+(!D C !B A)+(!D C B !A)+(!D C B A)), LSE_LINE_FILE_ID=3, LSE_LCOL=13, LSE_RCOL=44, LSE_LLINE=32, LSE_RLINE=32 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(11[2:53])
    defparam I1.init = 16'b0000000011111111;
    
endmodule
//
// Verilog Description of module inverter_U276
//

module inverter_U276 (\notGate[749]_keep , \notGate[750] ) /* synthesis syn_module_defined=1 */ ;
    input \notGate[749]_keep ;
    output \notGate[750] ;
    
    wire \notGate[749]_keep  /* synthesis alspreserve=1 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(25[15:22])
    
    LUT4 I1 (.A(\notGate[749]_keep ), .B(\notGate[749]_keep ), .C(\notGate[749]_keep ), 
         .D(\notGate[749]_keep ), .Z(\notGate[750] )) /* synthesis syn_instantiated=1, lut_function=((!D !C !B !A)+(!D !C !B A)+(!D !C B !A)+(!D !C B A)+(!D C !B !A)+(!D C !B A)+(!D C B !A)+(!D C B A)), LSE_LINE_FILE_ID=3, LSE_LCOL=13, LSE_RCOL=44, LSE_LLINE=32, LSE_RLINE=32 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(11[2:53])
    defparam I1.init = 16'b0000000011111111;
    
endmodule
//
// Verilog Description of module inverter_U277
//

module inverter_U277 (\notGate[73]_keep , \notGate[74] ) /* synthesis syn_module_defined=1 */ ;
    input \notGate[73]_keep ;
    output \notGate[74] ;
    
    wire \notGate[73]_keep  /* synthesis alspreserve=1 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(25[15:22])
    
    LUT4 I1 (.A(\notGate[73]_keep ), .B(\notGate[73]_keep ), .C(\notGate[73]_keep ), 
         .D(\notGate[73]_keep ), .Z(\notGate[74] )) /* synthesis syn_instantiated=1, lut_function=((!D !C !B !A)+(!D !C !B A)+(!D !C B !A)+(!D !C B A)+(!D C !B !A)+(!D C !B A)+(!D C B !A)+(!D C B A)), LSE_LINE_FILE_ID=3, LSE_LCOL=13, LSE_RCOL=44, LSE_LLINE=32, LSE_RLINE=32 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(11[2:53])
    defparam I1.init = 16'b0000000011111111;
    
endmodule
//
// Verilog Description of module inverter_U278
//

module inverter_U278 (\notGate[748]_keep , \notGate[749] ) /* synthesis syn_module_defined=1 */ ;
    input \notGate[748]_keep ;
    output \notGate[749] ;
    
    wire \notGate[748]_keep  /* synthesis alspreserve=1 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(25[15:22])
    
    LUT4 I1 (.A(\notGate[748]_keep ), .B(\notGate[748]_keep ), .C(\notGate[748]_keep ), 
         .D(\notGate[748]_keep ), .Z(\notGate[749] )) /* synthesis syn_instantiated=1, lut_function=((!D !C !B !A)+(!D !C !B A)+(!D !C B !A)+(!D !C B A)+(!D C !B !A)+(!D C !B A)+(!D C B !A)+(!D C B A)), LSE_LINE_FILE_ID=3, LSE_LCOL=13, LSE_RCOL=44, LSE_LLINE=32, LSE_RLINE=32 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(11[2:53])
    defparam I1.init = 16'b0000000011111111;
    
endmodule
//
// Verilog Description of module inverter_U279
//

module inverter_U279 (\notGate[747]_keep , \notGate[748] ) /* synthesis syn_module_defined=1 */ ;
    input \notGate[747]_keep ;
    output \notGate[748] ;
    
    wire \notGate[747]_keep  /* synthesis alspreserve=1 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(25[15:22])
    
    LUT4 I1 (.A(\notGate[747]_keep ), .B(\notGate[747]_keep ), .C(\notGate[747]_keep ), 
         .D(\notGate[747]_keep ), .Z(\notGate[748] )) /* synthesis syn_instantiated=1, lut_function=((!D !C !B !A)+(!D !C !B A)+(!D !C B !A)+(!D !C B A)+(!D C !B !A)+(!D C !B A)+(!D C B !A)+(!D C B A)), LSE_LINE_FILE_ID=3, LSE_LCOL=13, LSE_RCOL=44, LSE_LLINE=32, LSE_RLINE=32 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(11[2:53])
    defparam I1.init = 16'b0000000011111111;
    
endmodule
//
// Verilog Description of module inverter_U280
//

module inverter_U280 (\notGate[746]_keep , \notGate[747] ) /* synthesis syn_module_defined=1 */ ;
    input \notGate[746]_keep ;
    output \notGate[747] ;
    
    wire \notGate[746]_keep  /* synthesis alspreserve=1 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(25[15:22])
    
    LUT4 I1 (.A(\notGate[746]_keep ), .B(\notGate[746]_keep ), .C(\notGate[746]_keep ), 
         .D(\notGate[746]_keep ), .Z(\notGate[747] )) /* synthesis syn_instantiated=1, lut_function=((!D !C !B !A)+(!D !C !B A)+(!D !C B !A)+(!D !C B A)+(!D C !B !A)+(!D C !B A)+(!D C B !A)+(!D C B A)), LSE_LINE_FILE_ID=3, LSE_LCOL=13, LSE_RCOL=44, LSE_LLINE=32, LSE_RLINE=32 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(11[2:53])
    defparam I1.init = 16'b0000000011111111;
    
endmodule
//
// Verilog Description of module inverter_U281
//

module inverter_U281 (\notGate[745]_keep , \notGate[746] ) /* synthesis syn_module_defined=1 */ ;
    input \notGate[745]_keep ;
    output \notGate[746] ;
    
    wire \notGate[745]_keep  /* synthesis alspreserve=1 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(25[15:22])
    
    LUT4 I1 (.A(\notGate[745]_keep ), .B(\notGate[745]_keep ), .C(\notGate[745]_keep ), 
         .D(\notGate[745]_keep ), .Z(\notGate[746] )) /* synthesis syn_instantiated=1, lut_function=((!D !C !B !A)+(!D !C !B A)+(!D !C B !A)+(!D !C B A)+(!D C !B !A)+(!D C !B A)+(!D C B !A)+(!D C B A)), LSE_LINE_FILE_ID=3, LSE_LCOL=13, LSE_RCOL=44, LSE_LLINE=32, LSE_RLINE=32 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(11[2:53])
    defparam I1.init = 16'b0000000011111111;
    
endmodule
//
// Verilog Description of module inverter_U282
//

module inverter_U282 (\notGate[744]_keep , \notGate[745] ) /* synthesis syn_module_defined=1 */ ;
    input \notGate[744]_keep ;
    output \notGate[745] ;
    
    wire \notGate[744]_keep  /* synthesis alspreserve=1 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(25[15:22])
    
    LUT4 I1 (.A(\notGate[744]_keep ), .B(\notGate[744]_keep ), .C(\notGate[744]_keep ), 
         .D(\notGate[744]_keep ), .Z(\notGate[745] )) /* synthesis syn_instantiated=1, lut_function=((!D !C !B !A)+(!D !C !B A)+(!D !C B !A)+(!D !C B A)+(!D C !B !A)+(!D C !B A)+(!D C B !A)+(!D C B A)), LSE_LINE_FILE_ID=3, LSE_LCOL=13, LSE_RCOL=44, LSE_LLINE=32, LSE_RLINE=32 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(11[2:53])
    defparam I1.init = 16'b0000000011111111;
    
endmodule
//
// Verilog Description of module inverter_U283
//

module inverter_U283 (\notGate[743]_keep , \notGate[744] ) /* synthesis syn_module_defined=1 */ ;
    input \notGate[743]_keep ;
    output \notGate[744] ;
    
    wire \notGate[743]_keep  /* synthesis alspreserve=1 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(25[15:22])
    
    LUT4 I1 (.A(\notGate[743]_keep ), .B(\notGate[743]_keep ), .C(\notGate[743]_keep ), 
         .D(\notGate[743]_keep ), .Z(\notGate[744] )) /* synthesis syn_instantiated=1, lut_function=((!D !C !B !A)+(!D !C !B A)+(!D !C B !A)+(!D !C B A)+(!D C !B !A)+(!D C !B A)+(!D C B !A)+(!D C B A)), LSE_LINE_FILE_ID=3, LSE_LCOL=13, LSE_RCOL=44, LSE_LLINE=32, LSE_RLINE=32 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(11[2:53])
    defparam I1.init = 16'b0000000011111111;
    
endmodule
//
// Verilog Description of module inverter_U284
//

module inverter_U284 (\notGate[742]_keep , \notGate[743] ) /* synthesis syn_module_defined=1 */ ;
    input \notGate[742]_keep ;
    output \notGate[743] ;
    
    wire \notGate[742]_keep  /* synthesis alspreserve=1 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(25[15:22])
    
    LUT4 I1 (.A(\notGate[742]_keep ), .B(\notGate[742]_keep ), .C(\notGate[742]_keep ), 
         .D(\notGate[742]_keep ), .Z(\notGate[743] )) /* synthesis syn_instantiated=1, lut_function=((!D !C !B !A)+(!D !C !B A)+(!D !C B !A)+(!D !C B A)+(!D C !B !A)+(!D C !B A)+(!D C B !A)+(!D C B A)), LSE_LINE_FILE_ID=3, LSE_LCOL=13, LSE_RCOL=44, LSE_LLINE=32, LSE_RLINE=32 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(11[2:53])
    defparam I1.init = 16'b0000000011111111;
    
endmodule
//
// Verilog Description of module inverter_U285
//

module inverter_U285 (\notGate[741]_keep , \notGate[742] ) /* synthesis syn_module_defined=1 */ ;
    input \notGate[741]_keep ;
    output \notGate[742] ;
    
    wire \notGate[741]_keep  /* synthesis alspreserve=1 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(25[15:22])
    
    LUT4 I1 (.A(\notGate[741]_keep ), .B(\notGate[741]_keep ), .C(\notGate[741]_keep ), 
         .D(\notGate[741]_keep ), .Z(\notGate[742] )) /* synthesis syn_instantiated=1, lut_function=((!D !C !B !A)+(!D !C !B A)+(!D !C B !A)+(!D !C B A)+(!D C !B !A)+(!D C !B A)+(!D C B !A)+(!D C B A)), LSE_LINE_FILE_ID=3, LSE_LCOL=13, LSE_RCOL=44, LSE_LLINE=32, LSE_RLINE=32 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(11[2:53])
    defparam I1.init = 16'b0000000011111111;
    
endmodule
//
// Verilog Description of module inverter_U286
//

module inverter_U286 (\notGate[740]_keep , \notGate[741] ) /* synthesis syn_module_defined=1 */ ;
    input \notGate[740]_keep ;
    output \notGate[741] ;
    
    wire \notGate[740]_keep  /* synthesis alspreserve=1 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(25[15:22])
    
    LUT4 I1 (.A(\notGate[740]_keep ), .B(\notGate[740]_keep ), .C(\notGate[740]_keep ), 
         .D(\notGate[740]_keep ), .Z(\notGate[741] )) /* synthesis syn_instantiated=1, lut_function=((!D !C !B !A)+(!D !C !B A)+(!D !C B !A)+(!D !C B A)+(!D C !B !A)+(!D C !B A)+(!D C B !A)+(!D C B A)), LSE_LINE_FILE_ID=3, LSE_LCOL=13, LSE_RCOL=44, LSE_LLINE=32, LSE_RLINE=32 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(11[2:53])
    defparam I1.init = 16'b0000000011111111;
    
endmodule
//
// Verilog Description of module inverter_U287
//

module inverter_U287 (\notGate[739]_keep , \notGate[740] ) /* synthesis syn_module_defined=1 */ ;
    input \notGate[739]_keep ;
    output \notGate[740] ;
    
    wire \notGate[739]_keep  /* synthesis alspreserve=1 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(25[15:22])
    
    LUT4 I1 (.A(\notGate[739]_keep ), .B(\notGate[739]_keep ), .C(\notGate[739]_keep ), 
         .D(\notGate[739]_keep ), .Z(\notGate[740] )) /* synthesis syn_instantiated=1, lut_function=((!D !C !B !A)+(!D !C !B A)+(!D !C B !A)+(!D !C B A)+(!D C !B !A)+(!D C !B A)+(!D C B !A)+(!D C B A)), LSE_LINE_FILE_ID=3, LSE_LCOL=13, LSE_RCOL=44, LSE_LLINE=32, LSE_RLINE=32 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(11[2:53])
    defparam I1.init = 16'b0000000011111111;
    
endmodule
//
// Verilog Description of module inverter_U288
//

module inverter_U288 (\notGate[72]_keep , \notGate[73] ) /* synthesis syn_module_defined=1 */ ;
    input \notGate[72]_keep ;
    output \notGate[73] ;
    
    wire \notGate[72]_keep  /* synthesis alspreserve=1 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(25[15:22])
    
    LUT4 I1 (.A(\notGate[72]_keep ), .B(\notGate[72]_keep ), .C(\notGate[72]_keep ), 
         .D(\notGate[72]_keep ), .Z(\notGate[73] )) /* synthesis syn_instantiated=1, lut_function=((!D !C !B !A)+(!D !C !B A)+(!D !C B !A)+(!D !C B A)+(!D C !B !A)+(!D C !B A)+(!D C B !A)+(!D C B A)), LSE_LINE_FILE_ID=3, LSE_LCOL=13, LSE_RCOL=44, LSE_LLINE=32, LSE_RLINE=32 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(11[2:53])
    defparam I1.init = 16'b0000000011111111;
    
endmodule
//
// Verilog Description of module inverter_U289
//

module inverter_U289 (\notGate[738]_keep , \notGate[739] ) /* synthesis syn_module_defined=1 */ ;
    input \notGate[738]_keep ;
    output \notGate[739] ;
    
    wire \notGate[738]_keep  /* synthesis alspreserve=1 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(25[15:22])
    
    LUT4 I1 (.A(\notGate[738]_keep ), .B(\notGate[738]_keep ), .C(\notGate[738]_keep ), 
         .D(\notGate[738]_keep ), .Z(\notGate[739] )) /* synthesis syn_instantiated=1, lut_function=((!D !C !B !A)+(!D !C !B A)+(!D !C B !A)+(!D !C B A)+(!D C !B !A)+(!D C !B A)+(!D C B !A)+(!D C B A)), LSE_LINE_FILE_ID=3, LSE_LCOL=13, LSE_RCOL=44, LSE_LLINE=32, LSE_RLINE=32 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(11[2:53])
    defparam I1.init = 16'b0000000011111111;
    
endmodule
//
// Verilog Description of module inverter_U290
//

module inverter_U290 (\notGate[737]_keep , \notGate[738] ) /* synthesis syn_module_defined=1 */ ;
    input \notGate[737]_keep ;
    output \notGate[738] ;
    
    wire \notGate[737]_keep  /* synthesis alspreserve=1 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(25[15:22])
    
    LUT4 I1 (.A(\notGate[737]_keep ), .B(\notGate[737]_keep ), .C(\notGate[737]_keep ), 
         .D(\notGate[737]_keep ), .Z(\notGate[738] )) /* synthesis syn_instantiated=1, lut_function=((!D !C !B !A)+(!D !C !B A)+(!D !C B !A)+(!D !C B A)+(!D C !B !A)+(!D C !B A)+(!D C B !A)+(!D C B A)), LSE_LINE_FILE_ID=3, LSE_LCOL=13, LSE_RCOL=44, LSE_LLINE=32, LSE_RLINE=32 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(11[2:53])
    defparam I1.init = 16'b0000000011111111;
    
endmodule
//
// Verilog Description of module inverter_U291
//

module inverter_U291 (\notGate[736]_keep , \notGate[737] ) /* synthesis syn_module_defined=1 */ ;
    input \notGate[736]_keep ;
    output \notGate[737] ;
    
    wire \notGate[736]_keep  /* synthesis alspreserve=1 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(25[15:22])
    
    LUT4 I1 (.A(\notGate[736]_keep ), .B(\notGate[736]_keep ), .C(\notGate[736]_keep ), 
         .D(\notGate[736]_keep ), .Z(\notGate[737] )) /* synthesis syn_instantiated=1, lut_function=((!D !C !B !A)+(!D !C !B A)+(!D !C B !A)+(!D !C B A)+(!D C !B !A)+(!D C !B A)+(!D C B !A)+(!D C B A)), LSE_LINE_FILE_ID=3, LSE_LCOL=13, LSE_RCOL=44, LSE_LLINE=32, LSE_RLINE=32 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(11[2:53])
    defparam I1.init = 16'b0000000011111111;
    
endmodule
//
// Verilog Description of module inverter_U292
//

module inverter_U292 (\notGate[735]_keep , \notGate[736] ) /* synthesis syn_module_defined=1 */ ;
    input \notGate[735]_keep ;
    output \notGate[736] ;
    
    wire \notGate[735]_keep  /* synthesis alspreserve=1 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(25[15:22])
    
    LUT4 I1 (.A(\notGate[735]_keep ), .B(\notGate[735]_keep ), .C(\notGate[735]_keep ), 
         .D(\notGate[735]_keep ), .Z(\notGate[736] )) /* synthesis syn_instantiated=1, lut_function=((!D !C !B !A)+(!D !C !B A)+(!D !C B !A)+(!D !C B A)+(!D C !B !A)+(!D C !B A)+(!D C B !A)+(!D C B A)), LSE_LINE_FILE_ID=3, LSE_LCOL=13, LSE_RCOL=44, LSE_LLINE=32, LSE_RLINE=32 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(11[2:53])
    defparam I1.init = 16'b0000000011111111;
    
endmodule
//
// Verilog Description of module inverter_U293
//

module inverter_U293 (\notGate[734]_keep , \notGate[735] ) /* synthesis syn_module_defined=1 */ ;
    input \notGate[734]_keep ;
    output \notGate[735] ;
    
    wire \notGate[734]_keep  /* synthesis alspreserve=1 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(25[15:22])
    
    LUT4 I1 (.A(\notGate[734]_keep ), .B(\notGate[734]_keep ), .C(\notGate[734]_keep ), 
         .D(\notGate[734]_keep ), .Z(\notGate[735] )) /* synthesis syn_instantiated=1, lut_function=((!D !C !B !A)+(!D !C !B A)+(!D !C B !A)+(!D !C B A)+(!D C !B !A)+(!D C !B A)+(!D C B !A)+(!D C B A)), LSE_LINE_FILE_ID=3, LSE_LCOL=13, LSE_RCOL=44, LSE_LLINE=32, LSE_RLINE=32 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(11[2:53])
    defparam I1.init = 16'b0000000011111111;
    
endmodule
//
// Verilog Description of module inverter_U294
//

module inverter_U294 (\notGate[733]_keep , \notGate[734] ) /* synthesis syn_module_defined=1 */ ;
    input \notGate[733]_keep ;
    output \notGate[734] ;
    
    wire \notGate[733]_keep  /* synthesis alspreserve=1 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(25[15:22])
    
    LUT4 I1 (.A(\notGate[733]_keep ), .B(\notGate[733]_keep ), .C(\notGate[733]_keep ), 
         .D(\notGate[733]_keep ), .Z(\notGate[734] )) /* synthesis syn_instantiated=1, lut_function=((!D !C !B !A)+(!D !C !B A)+(!D !C B !A)+(!D !C B A)+(!D C !B !A)+(!D C !B A)+(!D C B !A)+(!D C B A)), LSE_LINE_FILE_ID=3, LSE_LCOL=13, LSE_RCOL=44, LSE_LLINE=32, LSE_RLINE=32 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(11[2:53])
    defparam I1.init = 16'b0000000011111111;
    
endmodule
//
// Verilog Description of module inverter_U295
//

module inverter_U295 (\notGate[732]_keep , \notGate[733] ) /* synthesis syn_module_defined=1 */ ;
    input \notGate[732]_keep ;
    output \notGate[733] ;
    
    wire \notGate[732]_keep  /* synthesis alspreserve=1 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(25[15:22])
    
    LUT4 I1 (.A(\notGate[732]_keep ), .B(\notGate[732]_keep ), .C(\notGate[732]_keep ), 
         .D(\notGate[732]_keep ), .Z(\notGate[733] )) /* synthesis syn_instantiated=1, lut_function=((!D !C !B !A)+(!D !C !B A)+(!D !C B !A)+(!D !C B A)+(!D C !B !A)+(!D C !B A)+(!D C B !A)+(!D C B A)), LSE_LINE_FILE_ID=3, LSE_LCOL=13, LSE_RCOL=44, LSE_LLINE=32, LSE_RLINE=32 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(11[2:53])
    defparam I1.init = 16'b0000000011111111;
    
endmodule
//
// Verilog Description of module inverter_U296
//

module inverter_U296 (\notGate[731]_keep , \notGate[732] ) /* synthesis syn_module_defined=1 */ ;
    input \notGate[731]_keep ;
    output \notGate[732] ;
    
    wire \notGate[731]_keep  /* synthesis alspreserve=1 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(25[15:22])
    
    LUT4 I1 (.A(\notGate[731]_keep ), .B(\notGate[731]_keep ), .C(\notGate[731]_keep ), 
         .D(\notGate[731]_keep ), .Z(\notGate[732] )) /* synthesis syn_instantiated=1, lut_function=((!D !C !B !A)+(!D !C !B A)+(!D !C B !A)+(!D !C B A)+(!D C !B !A)+(!D C !B A)+(!D C B !A)+(!D C B A)), LSE_LINE_FILE_ID=3, LSE_LCOL=13, LSE_RCOL=44, LSE_LLINE=32, LSE_RLINE=32 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(11[2:53])
    defparam I1.init = 16'b0000000011111111;
    
endmodule
//
// Verilog Description of module inverter_U297
//

module inverter_U297 (\notGate[730]_keep , \notGate[731] ) /* synthesis syn_module_defined=1 */ ;
    input \notGate[730]_keep ;
    output \notGate[731] ;
    
    wire \notGate[730]_keep  /* synthesis alspreserve=1 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(25[15:22])
    
    LUT4 I1 (.A(\notGate[730]_keep ), .B(\notGate[730]_keep ), .C(\notGate[730]_keep ), 
         .D(\notGate[730]_keep ), .Z(\notGate[731] )) /* synthesis syn_instantiated=1, lut_function=((!D !C !B !A)+(!D !C !B A)+(!D !C B !A)+(!D !C B A)+(!D C !B !A)+(!D C !B A)+(!D C B !A)+(!D C B A)), LSE_LINE_FILE_ID=3, LSE_LCOL=13, LSE_RCOL=44, LSE_LLINE=32, LSE_RLINE=32 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(11[2:53])
    defparam I1.init = 16'b0000000011111111;
    
endmodule
//
// Verilog Description of module inverter_U298
//

module inverter_U298 (\notGate[729]_keep , \notGate[730] ) /* synthesis syn_module_defined=1 */ ;
    input \notGate[729]_keep ;
    output \notGate[730] ;
    
    wire \notGate[729]_keep  /* synthesis alspreserve=1 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(25[15:22])
    
    LUT4 I1 (.A(\notGate[729]_keep ), .B(\notGate[729]_keep ), .C(\notGate[729]_keep ), 
         .D(\notGate[729]_keep ), .Z(\notGate[730] )) /* synthesis syn_instantiated=1, lut_function=((!D !C !B !A)+(!D !C !B A)+(!D !C B !A)+(!D !C B A)+(!D C !B !A)+(!D C !B A)+(!D C B !A)+(!D C B A)), LSE_LINE_FILE_ID=3, LSE_LCOL=13, LSE_RCOL=44, LSE_LLINE=32, LSE_RLINE=32 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(11[2:53])
    defparam I1.init = 16'b0000000011111111;
    
endmodule
//
// Verilog Description of module inverter_U299
//

module inverter_U299 (\notGate[71]_keep , \notGate[72] ) /* synthesis syn_module_defined=1 */ ;
    input \notGate[71]_keep ;
    output \notGate[72] ;
    
    wire \notGate[71]_keep  /* synthesis alspreserve=1 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(25[15:22])
    
    LUT4 I1 (.A(\notGate[71]_keep ), .B(\notGate[71]_keep ), .C(\notGate[71]_keep ), 
         .D(\notGate[71]_keep ), .Z(\notGate[72] )) /* synthesis syn_instantiated=1, lut_function=((!D !C !B !A)+(!D !C !B A)+(!D !C B !A)+(!D !C B A)+(!D C !B !A)+(!D C !B A)+(!D C B !A)+(!D C B A)), LSE_LINE_FILE_ID=3, LSE_LCOL=13, LSE_RCOL=44, LSE_LLINE=32, LSE_RLINE=32 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(11[2:53])
    defparam I1.init = 16'b0000000011111111;
    
endmodule
//
// Verilog Description of module inverter_U300
//

module inverter_U300 (\notGate[728]_keep , \notGate[729] ) /* synthesis syn_module_defined=1 */ ;
    input \notGate[728]_keep ;
    output \notGate[729] ;
    
    wire \notGate[728]_keep  /* synthesis alspreserve=1 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(25[15:22])
    
    LUT4 I1 (.A(\notGate[728]_keep ), .B(\notGate[728]_keep ), .C(\notGate[728]_keep ), 
         .D(\notGate[728]_keep ), .Z(\notGate[729] )) /* synthesis syn_instantiated=1, lut_function=((!D !C !B !A)+(!D !C !B A)+(!D !C B !A)+(!D !C B A)+(!D C !B !A)+(!D C !B A)+(!D C B !A)+(!D C B A)), LSE_LINE_FILE_ID=3, LSE_LCOL=13, LSE_RCOL=44, LSE_LLINE=32, LSE_RLINE=32 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(11[2:53])
    defparam I1.init = 16'b0000000011111111;
    
endmodule
//
// Verilog Description of module inverter_U301
//

module inverter_U301 (\notGate[727]_keep , \notGate[728] ) /* synthesis syn_module_defined=1 */ ;
    input \notGate[727]_keep ;
    output \notGate[728] ;
    
    wire \notGate[727]_keep  /* synthesis alspreserve=1 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(25[15:22])
    
    LUT4 I1 (.A(\notGate[727]_keep ), .B(\notGate[727]_keep ), .C(\notGate[727]_keep ), 
         .D(\notGate[727]_keep ), .Z(\notGate[728] )) /* synthesis syn_instantiated=1, lut_function=((!D !C !B !A)+(!D !C !B A)+(!D !C B !A)+(!D !C B A)+(!D C !B !A)+(!D C !B A)+(!D C B !A)+(!D C B A)), LSE_LINE_FILE_ID=3, LSE_LCOL=13, LSE_RCOL=44, LSE_LLINE=32, LSE_RLINE=32 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(11[2:53])
    defparam I1.init = 16'b0000000011111111;
    
endmodule
//
// Verilog Description of module inverter_U302
//

module inverter_U302 (\notGate[726]_keep , \notGate[727] ) /* synthesis syn_module_defined=1 */ ;
    input \notGate[726]_keep ;
    output \notGate[727] ;
    
    wire \notGate[726]_keep  /* synthesis alspreserve=1 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(25[15:22])
    
    LUT4 I1 (.A(\notGate[726]_keep ), .B(\notGate[726]_keep ), .C(\notGate[726]_keep ), 
         .D(\notGate[726]_keep ), .Z(\notGate[727] )) /* synthesis syn_instantiated=1, lut_function=((!D !C !B !A)+(!D !C !B A)+(!D !C B !A)+(!D !C B A)+(!D C !B !A)+(!D C !B A)+(!D C B !A)+(!D C B A)), LSE_LINE_FILE_ID=3, LSE_LCOL=13, LSE_RCOL=44, LSE_LLINE=32, LSE_RLINE=32 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(11[2:53])
    defparam I1.init = 16'b0000000011111111;
    
endmodule
//
// Verilog Description of module inverter_U303
//

module inverter_U303 (\notGate[725]_keep , \notGate[726] ) /* synthesis syn_module_defined=1 */ ;
    input \notGate[725]_keep ;
    output \notGate[726] ;
    
    wire \notGate[725]_keep  /* synthesis alspreserve=1 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(25[15:22])
    
    LUT4 I1 (.A(\notGate[725]_keep ), .B(\notGate[725]_keep ), .C(\notGate[725]_keep ), 
         .D(\notGate[725]_keep ), .Z(\notGate[726] )) /* synthesis syn_instantiated=1, lut_function=((!D !C !B !A)+(!D !C !B A)+(!D !C B !A)+(!D !C B A)+(!D C !B !A)+(!D C !B A)+(!D C B !A)+(!D C B A)), LSE_LINE_FILE_ID=3, LSE_LCOL=13, LSE_RCOL=44, LSE_LLINE=32, LSE_RLINE=32 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(11[2:53])
    defparam I1.init = 16'b0000000011111111;
    
endmodule
//
// Verilog Description of module inverter_U304
//

module inverter_U304 (\notGate[724]_keep , \notGate[725] ) /* synthesis syn_module_defined=1 */ ;
    input \notGate[724]_keep ;
    output \notGate[725] ;
    
    wire \notGate[724]_keep  /* synthesis alspreserve=1 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(25[15:22])
    
    LUT4 I1 (.A(\notGate[724]_keep ), .B(\notGate[724]_keep ), .C(\notGate[724]_keep ), 
         .D(\notGate[724]_keep ), .Z(\notGate[725] )) /* synthesis syn_instantiated=1, lut_function=((!D !C !B !A)+(!D !C !B A)+(!D !C B !A)+(!D !C B A)+(!D C !B !A)+(!D C !B A)+(!D C B !A)+(!D C B A)), LSE_LINE_FILE_ID=3, LSE_LCOL=13, LSE_RCOL=44, LSE_LLINE=32, LSE_RLINE=32 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(11[2:53])
    defparam I1.init = 16'b0000000011111111;
    
endmodule
//
// Verilog Description of module inverter_U305
//

module inverter_U305 (\notGate[723]_keep , \notGate[724] ) /* synthesis syn_module_defined=1 */ ;
    input \notGate[723]_keep ;
    output \notGate[724] ;
    
    wire \notGate[723]_keep  /* synthesis alspreserve=1 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(25[15:22])
    
    LUT4 I1 (.A(\notGate[723]_keep ), .B(\notGate[723]_keep ), .C(\notGate[723]_keep ), 
         .D(\notGate[723]_keep ), .Z(\notGate[724] )) /* synthesis syn_instantiated=1, lut_function=((!D !C !B !A)+(!D !C !B A)+(!D !C B !A)+(!D !C B A)+(!D C !B !A)+(!D C !B A)+(!D C B !A)+(!D C B A)), LSE_LINE_FILE_ID=3, LSE_LCOL=13, LSE_RCOL=44, LSE_LLINE=32, LSE_RLINE=32 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(11[2:53])
    defparam I1.init = 16'b0000000011111111;
    
endmodule
//
// Verilog Description of module inverter_U306
//

module inverter_U306 (\notGate[722]_keep , \notGate[723] ) /* synthesis syn_module_defined=1 */ ;
    input \notGate[722]_keep ;
    output \notGate[723] ;
    
    wire \notGate[722]_keep  /* synthesis alspreserve=1 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(25[15:22])
    
    LUT4 I1 (.A(\notGate[722]_keep ), .B(\notGate[722]_keep ), .C(\notGate[722]_keep ), 
         .D(\notGate[722]_keep ), .Z(\notGate[723] )) /* synthesis syn_instantiated=1, lut_function=((!D !C !B !A)+(!D !C !B A)+(!D !C B !A)+(!D !C B A)+(!D C !B !A)+(!D C !B A)+(!D C B !A)+(!D C B A)), LSE_LINE_FILE_ID=3, LSE_LCOL=13, LSE_RCOL=44, LSE_LLINE=32, LSE_RLINE=32 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(11[2:53])
    defparam I1.init = 16'b0000000011111111;
    
endmodule
//
// Verilog Description of module inverter_U307
//

module inverter_U307 (\notGate[721]_keep , \notGate[722] ) /* synthesis syn_module_defined=1 */ ;
    input \notGate[721]_keep ;
    output \notGate[722] ;
    
    wire \notGate[721]_keep  /* synthesis alspreserve=1 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(25[15:22])
    
    LUT4 I1 (.A(\notGate[721]_keep ), .B(\notGate[721]_keep ), .C(\notGate[721]_keep ), 
         .D(\notGate[721]_keep ), .Z(\notGate[722] )) /* synthesis syn_instantiated=1, lut_function=((!D !C !B !A)+(!D !C !B A)+(!D !C B !A)+(!D !C B A)+(!D C !B !A)+(!D C !B A)+(!D C B !A)+(!D C B A)), LSE_LINE_FILE_ID=3, LSE_LCOL=13, LSE_RCOL=44, LSE_LLINE=32, LSE_RLINE=32 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(11[2:53])
    defparam I1.init = 16'b0000000011111111;
    
endmodule
//
// Verilog Description of module inverter_U308
//

module inverter_U308 (\notGate[720]_keep , \notGate[721] ) /* synthesis syn_module_defined=1 */ ;
    input \notGate[720]_keep ;
    output \notGate[721] ;
    
    wire \notGate[720]_keep  /* synthesis alspreserve=1 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(25[15:22])
    
    LUT4 I1 (.A(\notGate[720]_keep ), .B(\notGate[720]_keep ), .C(\notGate[720]_keep ), 
         .D(\notGate[720]_keep ), .Z(\notGate[721] )) /* synthesis syn_instantiated=1, lut_function=((!D !C !B !A)+(!D !C !B A)+(!D !C B !A)+(!D !C B A)+(!D C !B !A)+(!D C !B A)+(!D C B !A)+(!D C B A)), LSE_LINE_FILE_ID=3, LSE_LCOL=13, LSE_RCOL=44, LSE_LLINE=32, LSE_RLINE=32 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(11[2:53])
    defparam I1.init = 16'b0000000011111111;
    
endmodule
//
// Verilog Description of module inverter_U309
//

module inverter_U309 (\notGate[719]_keep , \notGate[720] ) /* synthesis syn_module_defined=1 */ ;
    input \notGate[719]_keep ;
    output \notGate[720] ;
    
    wire \notGate[719]_keep  /* synthesis alspreserve=1 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(25[15:22])
    
    LUT4 I1 (.A(\notGate[719]_keep ), .B(\notGate[719]_keep ), .C(\notGate[719]_keep ), 
         .D(\notGate[719]_keep ), .Z(\notGate[720] )) /* synthesis syn_instantiated=1, lut_function=((!D !C !B !A)+(!D !C !B A)+(!D !C B !A)+(!D !C B A)+(!D C !B !A)+(!D C !B A)+(!D C B !A)+(!D C B A)), LSE_LINE_FILE_ID=3, LSE_LCOL=13, LSE_RCOL=44, LSE_LLINE=32, LSE_RLINE=32 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(11[2:53])
    defparam I1.init = 16'b0000000011111111;
    
endmodule
//
// Verilog Description of module inverter_U310
//

module inverter_U310 (\notGate[70]_keep , \notGate[71] ) /* synthesis syn_module_defined=1 */ ;
    input \notGate[70]_keep ;
    output \notGate[71] ;
    
    wire \notGate[70]_keep  /* synthesis alspreserve=1 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(25[15:22])
    
    LUT4 I1 (.A(\notGate[70]_keep ), .B(\notGate[70]_keep ), .C(\notGate[70]_keep ), 
         .D(\notGate[70]_keep ), .Z(\notGate[71] )) /* synthesis syn_instantiated=1, lut_function=((!D !C !B !A)+(!D !C !B A)+(!D !C B !A)+(!D !C B A)+(!D C !B !A)+(!D C !B A)+(!D C B !A)+(!D C B A)), LSE_LINE_FILE_ID=3, LSE_LCOL=13, LSE_RCOL=44, LSE_LLINE=32, LSE_RLINE=32 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(11[2:53])
    defparam I1.init = 16'b0000000011111111;
    
endmodule
//
// Verilog Description of module inverter_U311
//

module inverter_U311 (\notGate[718]_keep , \notGate[719] ) /* synthesis syn_module_defined=1 */ ;
    input \notGate[718]_keep ;
    output \notGate[719] ;
    
    wire \notGate[718]_keep  /* synthesis alspreserve=1 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(25[15:22])
    
    LUT4 I1 (.A(\notGate[718]_keep ), .B(\notGate[718]_keep ), .C(\notGate[718]_keep ), 
         .D(\notGate[718]_keep ), .Z(\notGate[719] )) /* synthesis syn_instantiated=1, lut_function=((!D !C !B !A)+(!D !C !B A)+(!D !C B !A)+(!D !C B A)+(!D C !B !A)+(!D C !B A)+(!D C B !A)+(!D C B A)), LSE_LINE_FILE_ID=3, LSE_LCOL=13, LSE_RCOL=44, LSE_LLINE=32, LSE_RLINE=32 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(11[2:53])
    defparam I1.init = 16'b0000000011111111;
    
endmodule
//
// Verilog Description of module inverter_U312
//

module inverter_U312 (\notGate[717]_keep , \notGate[718] ) /* synthesis syn_module_defined=1 */ ;
    input \notGate[717]_keep ;
    output \notGate[718] ;
    
    wire \notGate[717]_keep  /* synthesis alspreserve=1 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(25[15:22])
    
    LUT4 I1 (.A(\notGate[717]_keep ), .B(\notGate[717]_keep ), .C(\notGate[717]_keep ), 
         .D(\notGate[717]_keep ), .Z(\notGate[718] )) /* synthesis syn_instantiated=1, lut_function=((!D !C !B !A)+(!D !C !B A)+(!D !C B !A)+(!D !C B A)+(!D C !B !A)+(!D C !B A)+(!D C B !A)+(!D C B A)), LSE_LINE_FILE_ID=3, LSE_LCOL=13, LSE_RCOL=44, LSE_LLINE=32, LSE_RLINE=32 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(11[2:53])
    defparam I1.init = 16'b0000000011111111;
    
endmodule
//
// Verilog Description of module inverter_U313
//

module inverter_U313 (\notGate[716]_keep , \notGate[717] ) /* synthesis syn_module_defined=1 */ ;
    input \notGate[716]_keep ;
    output \notGate[717] ;
    
    wire \notGate[716]_keep  /* synthesis alspreserve=1 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(25[15:22])
    
    LUT4 I1 (.A(\notGate[716]_keep ), .B(\notGate[716]_keep ), .C(\notGate[716]_keep ), 
         .D(\notGate[716]_keep ), .Z(\notGate[717] )) /* synthesis syn_instantiated=1, lut_function=((!D !C !B !A)+(!D !C !B A)+(!D !C B !A)+(!D !C B A)+(!D C !B !A)+(!D C !B A)+(!D C B !A)+(!D C B A)), LSE_LINE_FILE_ID=3, LSE_LCOL=13, LSE_RCOL=44, LSE_LLINE=32, LSE_RLINE=32 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(11[2:53])
    defparam I1.init = 16'b0000000011111111;
    
endmodule
//
// Verilog Description of module inverter_U314
//

module inverter_U314 (\notGate[715]_keep , \notGate[716] ) /* synthesis syn_module_defined=1 */ ;
    input \notGate[715]_keep ;
    output \notGate[716] ;
    
    wire \notGate[715]_keep  /* synthesis alspreserve=1 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(25[15:22])
    
    LUT4 I1 (.A(\notGate[715]_keep ), .B(\notGate[715]_keep ), .C(\notGate[715]_keep ), 
         .D(\notGate[715]_keep ), .Z(\notGate[716] )) /* synthesis syn_instantiated=1, lut_function=((!D !C !B !A)+(!D !C !B A)+(!D !C B !A)+(!D !C B A)+(!D C !B !A)+(!D C !B A)+(!D C B !A)+(!D C B A)), LSE_LINE_FILE_ID=3, LSE_LCOL=13, LSE_RCOL=44, LSE_LLINE=32, LSE_RLINE=32 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(11[2:53])
    defparam I1.init = 16'b0000000011111111;
    
endmodule
//
// Verilog Description of module inverter_U315
//

module inverter_U315 (\notGate[714]_keep , \notGate[715] ) /* synthesis syn_module_defined=1 */ ;
    input \notGate[714]_keep ;
    output \notGate[715] ;
    
    wire \notGate[714]_keep  /* synthesis alspreserve=1 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(25[15:22])
    
    LUT4 I1 (.A(\notGate[714]_keep ), .B(\notGate[714]_keep ), .C(\notGate[714]_keep ), 
         .D(\notGate[714]_keep ), .Z(\notGate[715] )) /* synthesis syn_instantiated=1, lut_function=((!D !C !B !A)+(!D !C !B A)+(!D !C B !A)+(!D !C B A)+(!D C !B !A)+(!D C !B A)+(!D C B !A)+(!D C B A)), LSE_LINE_FILE_ID=3, LSE_LCOL=13, LSE_RCOL=44, LSE_LLINE=32, LSE_RLINE=32 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(11[2:53])
    defparam I1.init = 16'b0000000011111111;
    
endmodule
//
// Verilog Description of module inverter_U316
//

module inverter_U316 (\notGate[713]_keep , \notGate[714] ) /* synthesis syn_module_defined=1 */ ;
    input \notGate[713]_keep ;
    output \notGate[714] ;
    
    wire \notGate[713]_keep  /* synthesis alspreserve=1 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(25[15:22])
    
    LUT4 I1 (.A(\notGate[713]_keep ), .B(\notGate[713]_keep ), .C(\notGate[713]_keep ), 
         .D(\notGate[713]_keep ), .Z(\notGate[714] )) /* synthesis syn_instantiated=1, lut_function=((!D !C !B !A)+(!D !C !B A)+(!D !C B !A)+(!D !C B A)+(!D C !B !A)+(!D C !B A)+(!D C B !A)+(!D C B A)), LSE_LINE_FILE_ID=3, LSE_LCOL=13, LSE_RCOL=44, LSE_LLINE=32, LSE_RLINE=32 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(11[2:53])
    defparam I1.init = 16'b0000000011111111;
    
endmodule
//
// Verilog Description of module inverter_U317
//

module inverter_U317 (\notGate[712]_keep , \notGate[713] ) /* synthesis syn_module_defined=1 */ ;
    input \notGate[712]_keep ;
    output \notGate[713] ;
    
    wire \notGate[712]_keep  /* synthesis alspreserve=1 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(25[15:22])
    
    LUT4 I1 (.A(\notGate[712]_keep ), .B(\notGate[712]_keep ), .C(\notGate[712]_keep ), 
         .D(\notGate[712]_keep ), .Z(\notGate[713] )) /* synthesis syn_instantiated=1, lut_function=((!D !C !B !A)+(!D !C !B A)+(!D !C B !A)+(!D !C B A)+(!D C !B !A)+(!D C !B A)+(!D C B !A)+(!D C B A)), LSE_LINE_FILE_ID=3, LSE_LCOL=13, LSE_RCOL=44, LSE_LLINE=32, LSE_RLINE=32 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(11[2:53])
    defparam I1.init = 16'b0000000011111111;
    
endmodule
//
// Verilog Description of module inverter_U318
//

module inverter_U318 (\notGate[711]_keep , \notGate[712] ) /* synthesis syn_module_defined=1 */ ;
    input \notGate[711]_keep ;
    output \notGate[712] ;
    
    wire \notGate[711]_keep  /* synthesis alspreserve=1 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(25[15:22])
    
    LUT4 I1 (.A(\notGate[711]_keep ), .B(\notGate[711]_keep ), .C(\notGate[711]_keep ), 
         .D(\notGate[711]_keep ), .Z(\notGate[712] )) /* synthesis syn_instantiated=1, lut_function=((!D !C !B !A)+(!D !C !B A)+(!D !C B !A)+(!D !C B A)+(!D C !B !A)+(!D C !B A)+(!D C B !A)+(!D C B A)), LSE_LINE_FILE_ID=3, LSE_LCOL=13, LSE_RCOL=44, LSE_LLINE=32, LSE_RLINE=32 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(11[2:53])
    defparam I1.init = 16'b0000000011111111;
    
endmodule
//
// Verilog Description of module inverter_U319
//

module inverter_U319 (\notGate[710]_keep , \notGate[711] ) /* synthesis syn_module_defined=1 */ ;
    input \notGate[710]_keep ;
    output \notGate[711] ;
    
    wire \notGate[710]_keep  /* synthesis alspreserve=1 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(25[15:22])
    
    LUT4 I1 (.A(\notGate[710]_keep ), .B(\notGate[710]_keep ), .C(\notGate[710]_keep ), 
         .D(\notGate[710]_keep ), .Z(\notGate[711] )) /* synthesis syn_instantiated=1, lut_function=((!D !C !B !A)+(!D !C !B A)+(!D !C B !A)+(!D !C B A)+(!D C !B !A)+(!D C !B A)+(!D C B !A)+(!D C B A)), LSE_LINE_FILE_ID=3, LSE_LCOL=13, LSE_RCOL=44, LSE_LLINE=32, LSE_RLINE=32 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(11[2:53])
    defparam I1.init = 16'b0000000011111111;
    
endmodule
//
// Verilog Description of module inverter_U320
//

module inverter_U320 (\notGate[709]_keep , \notGate[710] ) /* synthesis syn_module_defined=1 */ ;
    input \notGate[709]_keep ;
    output \notGate[710] ;
    
    wire \notGate[709]_keep  /* synthesis alspreserve=1 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(25[15:22])
    
    LUT4 I1 (.A(\notGate[709]_keep ), .B(\notGate[709]_keep ), .C(\notGate[709]_keep ), 
         .D(\notGate[709]_keep ), .Z(\notGate[710] )) /* synthesis syn_instantiated=1, lut_function=((!D !C !B !A)+(!D !C !B A)+(!D !C B !A)+(!D !C B A)+(!D C !B !A)+(!D C !B A)+(!D C B !A)+(!D C B A)), LSE_LINE_FILE_ID=3, LSE_LCOL=13, LSE_RCOL=44, LSE_LLINE=32, LSE_RLINE=32 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(11[2:53])
    defparam I1.init = 16'b0000000011111111;
    
endmodule
//
// Verilog Description of module inverter_U321
//

module inverter_U321 (\notGate[69]_keep , \notGate[70] ) /* synthesis syn_module_defined=1 */ ;
    input \notGate[69]_keep ;
    output \notGate[70] ;
    
    wire \notGate[69]_keep  /* synthesis alspreserve=1 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(25[15:22])
    
    LUT4 I1 (.A(\notGate[69]_keep ), .B(\notGate[69]_keep ), .C(\notGate[69]_keep ), 
         .D(\notGate[69]_keep ), .Z(\notGate[70] )) /* synthesis syn_instantiated=1, lut_function=((!D !C !B !A)+(!D !C !B A)+(!D !C B !A)+(!D !C B A)+(!D C !B !A)+(!D C !B A)+(!D C B !A)+(!D C B A)), LSE_LINE_FILE_ID=3, LSE_LCOL=13, LSE_RCOL=44, LSE_LLINE=32, LSE_RLINE=32 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(11[2:53])
    defparam I1.init = 16'b0000000011111111;
    
endmodule
//
// Verilog Description of module inverter_U322
//

module inverter_U322 (\notGate[708]_keep , \notGate[709] ) /* synthesis syn_module_defined=1 */ ;
    input \notGate[708]_keep ;
    output \notGate[709] ;
    
    wire \notGate[708]_keep  /* synthesis alspreserve=1 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(25[15:22])
    
    LUT4 I1 (.A(\notGate[708]_keep ), .B(\notGate[708]_keep ), .C(\notGate[708]_keep ), 
         .D(\notGate[708]_keep ), .Z(\notGate[709] )) /* synthesis syn_instantiated=1, lut_function=((!D !C !B !A)+(!D !C !B A)+(!D !C B !A)+(!D !C B A)+(!D C !B !A)+(!D C !B A)+(!D C B !A)+(!D C B A)), LSE_LINE_FILE_ID=3, LSE_LCOL=13, LSE_RCOL=44, LSE_LLINE=32, LSE_RLINE=32 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(11[2:53])
    defparam I1.init = 16'b0000000011111111;
    
endmodule
//
// Verilog Description of module inverter_U323
//

module inverter_U323 (\notGate[707]_keep , \notGate[708] ) /* synthesis syn_module_defined=1 */ ;
    input \notGate[707]_keep ;
    output \notGate[708] ;
    
    wire \notGate[707]_keep  /* synthesis alspreserve=1 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(25[15:22])
    
    LUT4 I1 (.A(\notGate[707]_keep ), .B(\notGate[707]_keep ), .C(\notGate[707]_keep ), 
         .D(\notGate[707]_keep ), .Z(\notGate[708] )) /* synthesis syn_instantiated=1, lut_function=((!D !C !B !A)+(!D !C !B A)+(!D !C B !A)+(!D !C B A)+(!D C !B !A)+(!D C !B A)+(!D C B !A)+(!D C B A)), LSE_LINE_FILE_ID=3, LSE_LCOL=13, LSE_RCOL=44, LSE_LLINE=32, LSE_RLINE=32 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(11[2:53])
    defparam I1.init = 16'b0000000011111111;
    
endmodule
//
// Verilog Description of module inverter_U324
//

module inverter_U324 (\notGate[706]_keep , \notGate[707] ) /* synthesis syn_module_defined=1 */ ;
    input \notGate[706]_keep ;
    output \notGate[707] ;
    
    wire \notGate[706]_keep  /* synthesis alspreserve=1 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(25[15:22])
    
    LUT4 I1 (.A(\notGate[706]_keep ), .B(\notGate[706]_keep ), .C(\notGate[706]_keep ), 
         .D(\notGate[706]_keep ), .Z(\notGate[707] )) /* synthesis syn_instantiated=1, lut_function=((!D !C !B !A)+(!D !C !B A)+(!D !C B !A)+(!D !C B A)+(!D C !B !A)+(!D C !B A)+(!D C B !A)+(!D C B A)), LSE_LINE_FILE_ID=3, LSE_LCOL=13, LSE_RCOL=44, LSE_LLINE=32, LSE_RLINE=32 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(11[2:53])
    defparam I1.init = 16'b0000000011111111;
    
endmodule
//
// Verilog Description of module inverter_U325
//

module inverter_U325 (\notGate[705]_keep , \notGate[706] ) /* synthesis syn_module_defined=1 */ ;
    input \notGate[705]_keep ;
    output \notGate[706] ;
    
    wire \notGate[705]_keep  /* synthesis alspreserve=1 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(25[15:22])
    
    LUT4 I1 (.A(\notGate[705]_keep ), .B(\notGate[705]_keep ), .C(\notGate[705]_keep ), 
         .D(\notGate[705]_keep ), .Z(\notGate[706] )) /* synthesis syn_instantiated=1, lut_function=((!D !C !B !A)+(!D !C !B A)+(!D !C B !A)+(!D !C B A)+(!D C !B !A)+(!D C !B A)+(!D C B !A)+(!D C B A)), LSE_LINE_FILE_ID=3, LSE_LCOL=13, LSE_RCOL=44, LSE_LLINE=32, LSE_RLINE=32 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(11[2:53])
    defparam I1.init = 16'b0000000011111111;
    
endmodule
//
// Verilog Description of module inverter_U326
//

module inverter_U326 (\notGate[704]_keep , \notGate[705] ) /* synthesis syn_module_defined=1 */ ;
    input \notGate[704]_keep ;
    output \notGate[705] ;
    
    wire \notGate[704]_keep  /* synthesis alspreserve=1 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(25[15:22])
    
    LUT4 I1 (.A(\notGate[704]_keep ), .B(\notGate[704]_keep ), .C(\notGate[704]_keep ), 
         .D(\notGate[704]_keep ), .Z(\notGate[705] )) /* synthesis syn_instantiated=1, lut_function=((!D !C !B !A)+(!D !C !B A)+(!D !C B !A)+(!D !C B A)+(!D C !B !A)+(!D C !B A)+(!D C B !A)+(!D C B A)), LSE_LINE_FILE_ID=3, LSE_LCOL=13, LSE_RCOL=44, LSE_LLINE=32, LSE_RLINE=32 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(11[2:53])
    defparam I1.init = 16'b0000000011111111;
    
endmodule
//
// Verilog Description of module inverter_U327
//

module inverter_U327 (\notGate[703]_keep , \notGate[704] ) /* synthesis syn_module_defined=1 */ ;
    input \notGate[703]_keep ;
    output \notGate[704] ;
    
    wire \notGate[703]_keep  /* synthesis alspreserve=1 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(25[15:22])
    
    LUT4 I1 (.A(\notGate[703]_keep ), .B(\notGate[703]_keep ), .C(\notGate[703]_keep ), 
         .D(\notGate[703]_keep ), .Z(\notGate[704] )) /* synthesis syn_instantiated=1, lut_function=((!D !C !B !A)+(!D !C !B A)+(!D !C B !A)+(!D !C B A)+(!D C !B !A)+(!D C !B A)+(!D C B !A)+(!D C B A)), LSE_LINE_FILE_ID=3, LSE_LCOL=13, LSE_RCOL=44, LSE_LLINE=32, LSE_RLINE=32 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(11[2:53])
    defparam I1.init = 16'b0000000011111111;
    
endmodule
//
// Verilog Description of module inverter_U328
//

module inverter_U328 (\notGate[702]_keep , \notGate[703] ) /* synthesis syn_module_defined=1 */ ;
    input \notGate[702]_keep ;
    output \notGate[703] ;
    
    wire \notGate[702]_keep  /* synthesis alspreserve=1 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(25[15:22])
    
    LUT4 I1 (.A(\notGate[702]_keep ), .B(\notGate[702]_keep ), .C(\notGate[702]_keep ), 
         .D(\notGate[702]_keep ), .Z(\notGate[703] )) /* synthesis syn_instantiated=1, lut_function=((!D !C !B !A)+(!D !C !B A)+(!D !C B !A)+(!D !C B A)+(!D C !B !A)+(!D C !B A)+(!D C B !A)+(!D C B A)), LSE_LINE_FILE_ID=3, LSE_LCOL=13, LSE_RCOL=44, LSE_LLINE=32, LSE_RLINE=32 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(11[2:53])
    defparam I1.init = 16'b0000000011111111;
    
endmodule
//
// Verilog Description of module inverter_U329
//

module inverter_U329 (\notGate[701]_keep , \notGate[702] ) /* synthesis syn_module_defined=1 */ ;
    input \notGate[701]_keep ;
    output \notGate[702] ;
    
    wire \notGate[701]_keep  /* synthesis alspreserve=1 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(25[15:22])
    
    LUT4 I1 (.A(\notGate[701]_keep ), .B(\notGate[701]_keep ), .C(\notGate[701]_keep ), 
         .D(\notGate[701]_keep ), .Z(\notGate[702] )) /* synthesis syn_instantiated=1, lut_function=((!D !C !B !A)+(!D !C !B A)+(!D !C B !A)+(!D !C B A)+(!D C !B !A)+(!D C !B A)+(!D C B !A)+(!D C B A)), LSE_LINE_FILE_ID=3, LSE_LCOL=13, LSE_RCOL=44, LSE_LLINE=32, LSE_RLINE=32 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(11[2:53])
    defparam I1.init = 16'b0000000011111111;
    
endmodule
//
// Verilog Description of module inverter_U330
//

module inverter_U330 (\notGate[700]_keep , \notGate[701] ) /* synthesis syn_module_defined=1 */ ;
    input \notGate[700]_keep ;
    output \notGate[701] ;
    
    wire \notGate[700]_keep  /* synthesis alspreserve=1 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(25[15:22])
    
    LUT4 I1 (.A(\notGate[700]_keep ), .B(\notGate[700]_keep ), .C(\notGate[700]_keep ), 
         .D(\notGate[700]_keep ), .Z(\notGate[701] )) /* synthesis syn_instantiated=1, lut_function=((!D !C !B !A)+(!D !C !B A)+(!D !C B !A)+(!D !C B A)+(!D C !B !A)+(!D C !B A)+(!D C B !A)+(!D C B A)), LSE_LINE_FILE_ID=3, LSE_LCOL=13, LSE_RCOL=44, LSE_LLINE=32, LSE_RLINE=32 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(11[2:53])
    defparam I1.init = 16'b0000000011111111;
    
endmodule
//
// Verilog Description of module inverter_U331
//

module inverter_U331 (\notGate[699]_keep , \notGate[700] ) /* synthesis syn_module_defined=1 */ ;
    input \notGate[699]_keep ;
    output \notGate[700] ;
    
    wire \notGate[699]_keep  /* synthesis alspreserve=1 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(25[15:22])
    
    LUT4 I1 (.A(\notGate[699]_keep ), .B(\notGate[699]_keep ), .C(\notGate[699]_keep ), 
         .D(\notGate[699]_keep ), .Z(\notGate[700] )) /* synthesis syn_instantiated=1, lut_function=((!D !C !B !A)+(!D !C !B A)+(!D !C B !A)+(!D !C B A)+(!D C !B !A)+(!D C !B A)+(!D C B !A)+(!D C B A)), LSE_LINE_FILE_ID=3, LSE_LCOL=13, LSE_RCOL=44, LSE_LLINE=32, LSE_RLINE=32 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(11[2:53])
    defparam I1.init = 16'b0000000011111111;
    
endmodule
//
// Verilog Description of module inverter_U332
//

module inverter_U332 (\notGate[5]_keep , \notGate[6] ) /* synthesis syn_module_defined=1 */ ;
    input \notGate[5]_keep ;
    output \notGate[6] ;
    
    wire \notGate[5]_keep  /* synthesis alspreserve=1 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(25[15:22])
    
    LUT4 I1 (.A(\notGate[5]_keep ), .B(\notGate[5]_keep ), .C(\notGate[5]_keep ), 
         .D(\notGate[5]_keep ), .Z(\notGate[6] )) /* synthesis syn_instantiated=1, lut_function=((!D !C !B !A)+(!D !C !B A)+(!D !C B !A)+(!D !C B A)+(!D C !B !A)+(!D C !B A)+(!D C B !A)+(!D C B A)), LSE_LINE_FILE_ID=3, LSE_LCOL=13, LSE_RCOL=44, LSE_LLINE=32, LSE_RLINE=32 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(11[2:53])
    defparam I1.init = 16'b0000000011111111;
    
endmodule
//
// Verilog Description of module inverter_U333
//

module inverter_U333 (\notGate[68]_keep , \notGate[69] ) /* synthesis syn_module_defined=1 */ ;
    input \notGate[68]_keep ;
    output \notGate[69] ;
    
    wire \notGate[68]_keep  /* synthesis alspreserve=1 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(25[15:22])
    
    LUT4 I1 (.A(\notGate[68]_keep ), .B(\notGate[68]_keep ), .C(\notGate[68]_keep ), 
         .D(\notGate[68]_keep ), .Z(\notGate[69] )) /* synthesis syn_instantiated=1, lut_function=((!D !C !B !A)+(!D !C !B A)+(!D !C B !A)+(!D !C B A)+(!D C !B !A)+(!D C !B A)+(!D C B !A)+(!D C B A)), LSE_LINE_FILE_ID=3, LSE_LCOL=13, LSE_RCOL=44, LSE_LLINE=32, LSE_RLINE=32 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(11[2:53])
    defparam I1.init = 16'b0000000011111111;
    
endmodule
//
// Verilog Description of module inverter_U334
//

module inverter_U334 (\notGate[698]_keep , \notGate[699] ) /* synthesis syn_module_defined=1 */ ;
    input \notGate[698]_keep ;
    output \notGate[699] ;
    
    wire \notGate[698]_keep  /* synthesis alspreserve=1 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(25[15:22])
    
    LUT4 I1 (.A(\notGate[698]_keep ), .B(\notGate[698]_keep ), .C(\notGate[698]_keep ), 
         .D(\notGate[698]_keep ), .Z(\notGate[699] )) /* synthesis syn_instantiated=1, lut_function=((!D !C !B !A)+(!D !C !B A)+(!D !C B !A)+(!D !C B A)+(!D C !B !A)+(!D C !B A)+(!D C B !A)+(!D C B A)), LSE_LINE_FILE_ID=3, LSE_LCOL=13, LSE_RCOL=44, LSE_LLINE=32, LSE_RLINE=32 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(11[2:53])
    defparam I1.init = 16'b0000000011111111;
    
endmodule
//
// Verilog Description of module inverter_U335
//

module inverter_U335 (\notGate[697]_keep , \notGate[698] ) /* synthesis syn_module_defined=1 */ ;
    input \notGate[697]_keep ;
    output \notGate[698] ;
    
    wire \notGate[697]_keep  /* synthesis alspreserve=1 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(25[15:22])
    
    LUT4 I1 (.A(\notGate[697]_keep ), .B(\notGate[697]_keep ), .C(\notGate[697]_keep ), 
         .D(\notGate[697]_keep ), .Z(\notGate[698] )) /* synthesis syn_instantiated=1, lut_function=((!D !C !B !A)+(!D !C !B A)+(!D !C B !A)+(!D !C B A)+(!D C !B !A)+(!D C !B A)+(!D C B !A)+(!D C B A)), LSE_LINE_FILE_ID=3, LSE_LCOL=13, LSE_RCOL=44, LSE_LLINE=32, LSE_RLINE=32 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(11[2:53])
    defparam I1.init = 16'b0000000011111111;
    
endmodule
//
// Verilog Description of module inverter_U336
//

module inverter_U336 (\notGate[696]_keep , \notGate[697] ) /* synthesis syn_module_defined=1 */ ;
    input \notGate[696]_keep ;
    output \notGate[697] ;
    
    wire \notGate[696]_keep  /* synthesis alspreserve=1 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(25[15:22])
    
    LUT4 I1 (.A(\notGate[696]_keep ), .B(\notGate[696]_keep ), .C(\notGate[696]_keep ), 
         .D(\notGate[696]_keep ), .Z(\notGate[697] )) /* synthesis syn_instantiated=1, lut_function=((!D !C !B !A)+(!D !C !B A)+(!D !C B !A)+(!D !C B A)+(!D C !B !A)+(!D C !B A)+(!D C B !A)+(!D C B A)), LSE_LINE_FILE_ID=3, LSE_LCOL=13, LSE_RCOL=44, LSE_LLINE=32, LSE_RLINE=32 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(11[2:53])
    defparam I1.init = 16'b0000000011111111;
    
endmodule
//
// Verilog Description of module inverter_U337
//

module inverter_U337 (\notGate[695]_keep , \notGate[696] ) /* synthesis syn_module_defined=1 */ ;
    input \notGate[695]_keep ;
    output \notGate[696] ;
    
    wire \notGate[695]_keep  /* synthesis alspreserve=1 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(25[15:22])
    
    LUT4 I1 (.A(\notGate[695]_keep ), .B(\notGate[695]_keep ), .C(\notGate[695]_keep ), 
         .D(\notGate[695]_keep ), .Z(\notGate[696] )) /* synthesis syn_instantiated=1, lut_function=((!D !C !B !A)+(!D !C !B A)+(!D !C B !A)+(!D !C B A)+(!D C !B !A)+(!D C !B A)+(!D C B !A)+(!D C B A)), LSE_LINE_FILE_ID=3, LSE_LCOL=13, LSE_RCOL=44, LSE_LLINE=32, LSE_RLINE=32 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(11[2:53])
    defparam I1.init = 16'b0000000011111111;
    
endmodule
//
// Verilog Description of module inverter_U338
//

module inverter_U338 (\notGate[694]_keep , \notGate[695] ) /* synthesis syn_module_defined=1 */ ;
    input \notGate[694]_keep ;
    output \notGate[695] ;
    
    wire \notGate[694]_keep  /* synthesis alspreserve=1 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(25[15:22])
    
    LUT4 I1 (.A(\notGate[694]_keep ), .B(\notGate[694]_keep ), .C(\notGate[694]_keep ), 
         .D(\notGate[694]_keep ), .Z(\notGate[695] )) /* synthesis syn_instantiated=1, lut_function=((!D !C !B !A)+(!D !C !B A)+(!D !C B !A)+(!D !C B A)+(!D C !B !A)+(!D C !B A)+(!D C B !A)+(!D C B A)), LSE_LINE_FILE_ID=3, LSE_LCOL=13, LSE_RCOL=44, LSE_LLINE=32, LSE_RLINE=32 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(11[2:53])
    defparam I1.init = 16'b0000000011111111;
    
endmodule
//
// Verilog Description of module inverter_U339
//

module inverter_U339 (\notGate[693]_keep , \notGate[694] ) /* synthesis syn_module_defined=1 */ ;
    input \notGate[693]_keep ;
    output \notGate[694] ;
    
    wire \notGate[693]_keep  /* synthesis alspreserve=1 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(25[15:22])
    
    LUT4 I1 (.A(\notGate[693]_keep ), .B(\notGate[693]_keep ), .C(\notGate[693]_keep ), 
         .D(\notGate[693]_keep ), .Z(\notGate[694] )) /* synthesis syn_instantiated=1, lut_function=((!D !C !B !A)+(!D !C !B A)+(!D !C B !A)+(!D !C B A)+(!D C !B !A)+(!D C !B A)+(!D C B !A)+(!D C B A)), LSE_LINE_FILE_ID=3, LSE_LCOL=13, LSE_RCOL=44, LSE_LLINE=32, LSE_RLINE=32 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(11[2:53])
    defparam I1.init = 16'b0000000011111111;
    
endmodule
//
// Verilog Description of module inverter_U340
//

module inverter_U340 (\notGate[692]_keep , \notGate[693] ) /* synthesis syn_module_defined=1 */ ;
    input \notGate[692]_keep ;
    output \notGate[693] ;
    
    wire \notGate[692]_keep  /* synthesis alspreserve=1 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(25[15:22])
    
    LUT4 I1 (.A(\notGate[692]_keep ), .B(\notGate[692]_keep ), .C(\notGate[692]_keep ), 
         .D(\notGate[692]_keep ), .Z(\notGate[693] )) /* synthesis syn_instantiated=1, lut_function=((!D !C !B !A)+(!D !C !B A)+(!D !C B !A)+(!D !C B A)+(!D C !B !A)+(!D C !B A)+(!D C B !A)+(!D C B A)), LSE_LINE_FILE_ID=3, LSE_LCOL=13, LSE_RCOL=44, LSE_LLINE=32, LSE_RLINE=32 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(11[2:53])
    defparam I1.init = 16'b0000000011111111;
    
endmodule
//
// Verilog Description of module inverter_U341
//

module inverter_U341 (\notGate[691]_keep , \notGate[692] ) /* synthesis syn_module_defined=1 */ ;
    input \notGate[691]_keep ;
    output \notGate[692] ;
    
    wire \notGate[691]_keep  /* synthesis alspreserve=1 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(25[15:22])
    
    LUT4 I1 (.A(\notGate[691]_keep ), .B(\notGate[691]_keep ), .C(\notGate[691]_keep ), 
         .D(\notGate[691]_keep ), .Z(\notGate[692] )) /* synthesis syn_instantiated=1, lut_function=((!D !C !B !A)+(!D !C !B A)+(!D !C B !A)+(!D !C B A)+(!D C !B !A)+(!D C !B A)+(!D C B !A)+(!D C B A)), LSE_LINE_FILE_ID=3, LSE_LCOL=13, LSE_RCOL=44, LSE_LLINE=32, LSE_RLINE=32 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(11[2:53])
    defparam I1.init = 16'b0000000011111111;
    
endmodule
//
// Verilog Description of module inverter_U342
//

module inverter_U342 (\notGate[690]_keep , \notGate[691] ) /* synthesis syn_module_defined=1 */ ;
    input \notGate[690]_keep ;
    output \notGate[691] ;
    
    wire \notGate[690]_keep  /* synthesis alspreserve=1 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(25[15:22])
    
    LUT4 I1 (.A(\notGate[690]_keep ), .B(\notGate[690]_keep ), .C(\notGate[690]_keep ), 
         .D(\notGate[690]_keep ), .Z(\notGate[691] )) /* synthesis syn_instantiated=1, lut_function=((!D !C !B !A)+(!D !C !B A)+(!D !C B !A)+(!D !C B A)+(!D C !B !A)+(!D C !B A)+(!D C B !A)+(!D C B A)), LSE_LINE_FILE_ID=3, LSE_LCOL=13, LSE_RCOL=44, LSE_LLINE=32, LSE_RLINE=32 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(11[2:53])
    defparam I1.init = 16'b0000000011111111;
    
endmodule
//
// Verilog Description of module inverter_U343
//

module inverter_U343 (\notGate[689]_keep , \notGate[690] ) /* synthesis syn_module_defined=1 */ ;
    input \notGate[689]_keep ;
    output \notGate[690] ;
    
    wire \notGate[689]_keep  /* synthesis alspreserve=1 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(25[15:22])
    
    LUT4 I1 (.A(\notGate[689]_keep ), .B(\notGate[689]_keep ), .C(\notGate[689]_keep ), 
         .D(\notGate[689]_keep ), .Z(\notGate[690] )) /* synthesis syn_instantiated=1, lut_function=((!D !C !B !A)+(!D !C !B A)+(!D !C B !A)+(!D !C B A)+(!D C !B !A)+(!D C !B A)+(!D C B !A)+(!D C B A)), LSE_LINE_FILE_ID=3, LSE_LCOL=13, LSE_RCOL=44, LSE_LLINE=32, LSE_RLINE=32 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(11[2:53])
    defparam I1.init = 16'b0000000011111111;
    
endmodule
//
// Verilog Description of module inverter_U344
//

module inverter_U344 (\notGate[67]_keep , \notGate[68] ) /* synthesis syn_module_defined=1 */ ;
    input \notGate[67]_keep ;
    output \notGate[68] ;
    
    wire \notGate[67]_keep  /* synthesis alspreserve=1 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(25[15:22])
    
    LUT4 I1 (.A(\notGate[67]_keep ), .B(\notGate[67]_keep ), .C(\notGate[67]_keep ), 
         .D(\notGate[67]_keep ), .Z(\notGate[68] )) /* synthesis syn_instantiated=1, lut_function=((!D !C !B !A)+(!D !C !B A)+(!D !C B !A)+(!D !C B A)+(!D C !B !A)+(!D C !B A)+(!D C B !A)+(!D C B A)), LSE_LINE_FILE_ID=3, LSE_LCOL=13, LSE_RCOL=44, LSE_LLINE=32, LSE_RLINE=32 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(11[2:53])
    defparam I1.init = 16'b0000000011111111;
    
endmodule
//
// Verilog Description of module inverter_U345
//

module inverter_U345 (\notGate[688]_keep , \notGate[689] ) /* synthesis syn_module_defined=1 */ ;
    input \notGate[688]_keep ;
    output \notGate[689] ;
    
    wire \notGate[688]_keep  /* synthesis alspreserve=1 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(25[15:22])
    
    LUT4 I1 (.A(\notGate[688]_keep ), .B(\notGate[688]_keep ), .C(\notGate[688]_keep ), 
         .D(\notGate[688]_keep ), .Z(\notGate[689] )) /* synthesis syn_instantiated=1, lut_function=((!D !C !B !A)+(!D !C !B A)+(!D !C B !A)+(!D !C B A)+(!D C !B !A)+(!D C !B A)+(!D C B !A)+(!D C B A)), LSE_LINE_FILE_ID=3, LSE_LCOL=13, LSE_RCOL=44, LSE_LLINE=32, LSE_RLINE=32 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(11[2:53])
    defparam I1.init = 16'b0000000011111111;
    
endmodule
//
// Verilog Description of module inverter_U346
//

module inverter_U346 (\notGate[687]_keep , \notGate[688] ) /* synthesis syn_module_defined=1 */ ;
    input \notGate[687]_keep ;
    output \notGate[688] ;
    
    wire \notGate[687]_keep  /* synthesis alspreserve=1 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(25[15:22])
    
    LUT4 I1 (.A(\notGate[687]_keep ), .B(\notGate[687]_keep ), .C(\notGate[687]_keep ), 
         .D(\notGate[687]_keep ), .Z(\notGate[688] )) /* synthesis syn_instantiated=1, lut_function=((!D !C !B !A)+(!D !C !B A)+(!D !C B !A)+(!D !C B A)+(!D C !B !A)+(!D C !B A)+(!D C B !A)+(!D C B A)), LSE_LINE_FILE_ID=3, LSE_LCOL=13, LSE_RCOL=44, LSE_LLINE=32, LSE_RLINE=32 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(11[2:53])
    defparam I1.init = 16'b0000000011111111;
    
endmodule
//
// Verilog Description of module inverter_U347
//

module inverter_U347 (\notGate[686]_keep , \notGate[687] ) /* synthesis syn_module_defined=1 */ ;
    input \notGate[686]_keep ;
    output \notGate[687] ;
    
    wire \notGate[686]_keep  /* synthesis alspreserve=1 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(25[15:22])
    
    LUT4 I1 (.A(\notGate[686]_keep ), .B(\notGate[686]_keep ), .C(\notGate[686]_keep ), 
         .D(\notGate[686]_keep ), .Z(\notGate[687] )) /* synthesis syn_instantiated=1, lut_function=((!D !C !B !A)+(!D !C !B A)+(!D !C B !A)+(!D !C B A)+(!D C !B !A)+(!D C !B A)+(!D C B !A)+(!D C B A)), LSE_LINE_FILE_ID=3, LSE_LCOL=13, LSE_RCOL=44, LSE_LLINE=32, LSE_RLINE=32 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(11[2:53])
    defparam I1.init = 16'b0000000011111111;
    
endmodule
//
// Verilog Description of module inverter_U348
//

module inverter_U348 (\notGate[685]_keep , \notGate[686] ) /* synthesis syn_module_defined=1 */ ;
    input \notGate[685]_keep ;
    output \notGate[686] ;
    
    wire \notGate[685]_keep  /* synthesis alspreserve=1 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(25[15:22])
    
    LUT4 I1 (.A(\notGate[685]_keep ), .B(\notGate[685]_keep ), .C(\notGate[685]_keep ), 
         .D(\notGate[685]_keep ), .Z(\notGate[686] )) /* synthesis syn_instantiated=1, lut_function=((!D !C !B !A)+(!D !C !B A)+(!D !C B !A)+(!D !C B A)+(!D C !B !A)+(!D C !B A)+(!D C B !A)+(!D C B A)), LSE_LINE_FILE_ID=3, LSE_LCOL=13, LSE_RCOL=44, LSE_LLINE=32, LSE_RLINE=32 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(11[2:53])
    defparam I1.init = 16'b0000000011111111;
    
endmodule
//
// Verilog Description of module inverter_U349
//

module inverter_U349 (\notGate[684]_keep , \notGate[685] ) /* synthesis syn_module_defined=1 */ ;
    input \notGate[684]_keep ;
    output \notGate[685] ;
    
    wire \notGate[684]_keep  /* synthesis alspreserve=1 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(25[15:22])
    
    LUT4 I1 (.A(\notGate[684]_keep ), .B(\notGate[684]_keep ), .C(\notGate[684]_keep ), 
         .D(\notGate[684]_keep ), .Z(\notGate[685] )) /* synthesis syn_instantiated=1, lut_function=((!D !C !B !A)+(!D !C !B A)+(!D !C B !A)+(!D !C B A)+(!D C !B !A)+(!D C !B A)+(!D C B !A)+(!D C B A)), LSE_LINE_FILE_ID=3, LSE_LCOL=13, LSE_RCOL=44, LSE_LLINE=32, LSE_RLINE=32 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(11[2:53])
    defparam I1.init = 16'b0000000011111111;
    
endmodule
//
// Verilog Description of module inverter_U350
//

module inverter_U350 (\notGate[683]_keep , \notGate[684] ) /* synthesis syn_module_defined=1 */ ;
    input \notGate[683]_keep ;
    output \notGate[684] ;
    
    wire \notGate[683]_keep  /* synthesis alspreserve=1 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(25[15:22])
    
    LUT4 I1 (.A(\notGate[683]_keep ), .B(\notGate[683]_keep ), .C(\notGate[683]_keep ), 
         .D(\notGate[683]_keep ), .Z(\notGate[684] )) /* synthesis syn_instantiated=1, lut_function=((!D !C !B !A)+(!D !C !B A)+(!D !C B !A)+(!D !C B A)+(!D C !B !A)+(!D C !B A)+(!D C B !A)+(!D C B A)), LSE_LINE_FILE_ID=3, LSE_LCOL=13, LSE_RCOL=44, LSE_LLINE=32, LSE_RLINE=32 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(11[2:53])
    defparam I1.init = 16'b0000000011111111;
    
endmodule
//
// Verilog Description of module inverter_U351
//

module inverter_U351 (\notGate[682]_keep , \notGate[683] ) /* synthesis syn_module_defined=1 */ ;
    input \notGate[682]_keep ;
    output \notGate[683] ;
    
    wire \notGate[682]_keep  /* synthesis alspreserve=1 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(25[15:22])
    
    LUT4 I1 (.A(\notGate[682]_keep ), .B(\notGate[682]_keep ), .C(\notGate[682]_keep ), 
         .D(\notGate[682]_keep ), .Z(\notGate[683] )) /* synthesis syn_instantiated=1, lut_function=((!D !C !B !A)+(!D !C !B A)+(!D !C B !A)+(!D !C B A)+(!D C !B !A)+(!D C !B A)+(!D C B !A)+(!D C B A)), LSE_LINE_FILE_ID=3, LSE_LCOL=13, LSE_RCOL=44, LSE_LLINE=32, LSE_RLINE=32 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(11[2:53])
    defparam I1.init = 16'b0000000011111111;
    
endmodule
//
// Verilog Description of module inverter_U352
//

module inverter_U352 (\notGate[681]_keep , \notGate[682] ) /* synthesis syn_module_defined=1 */ ;
    input \notGate[681]_keep ;
    output \notGate[682] ;
    
    wire \notGate[681]_keep  /* synthesis alspreserve=1 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(25[15:22])
    
    LUT4 I1 (.A(\notGate[681]_keep ), .B(\notGate[681]_keep ), .C(\notGate[681]_keep ), 
         .D(\notGate[681]_keep ), .Z(\notGate[682] )) /* synthesis syn_instantiated=1, lut_function=((!D !C !B !A)+(!D !C !B A)+(!D !C B !A)+(!D !C B A)+(!D C !B !A)+(!D C !B A)+(!D C B !A)+(!D C B A)), LSE_LINE_FILE_ID=3, LSE_LCOL=13, LSE_RCOL=44, LSE_LLINE=32, LSE_RLINE=32 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(11[2:53])
    defparam I1.init = 16'b0000000011111111;
    
endmodule
//
// Verilog Description of module inverter_U353
//

module inverter_U353 (\notGate[680]_keep , \notGate[681] ) /* synthesis syn_module_defined=1 */ ;
    input \notGate[680]_keep ;
    output \notGate[681] ;
    
    wire \notGate[680]_keep  /* synthesis alspreserve=1 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(25[15:22])
    
    LUT4 I1 (.A(\notGate[680]_keep ), .B(\notGate[680]_keep ), .C(\notGate[680]_keep ), 
         .D(\notGate[680]_keep ), .Z(\notGate[681] )) /* synthesis syn_instantiated=1, lut_function=((!D !C !B !A)+(!D !C !B A)+(!D !C B !A)+(!D !C B A)+(!D C !B !A)+(!D C !B A)+(!D C B !A)+(!D C B A)), LSE_LINE_FILE_ID=3, LSE_LCOL=13, LSE_RCOL=44, LSE_LLINE=32, LSE_RLINE=32 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(11[2:53])
    defparam I1.init = 16'b0000000011111111;
    
endmodule
//
// Verilog Description of module inverter_U354
//

module inverter_U354 (\notGate[679]_keep , \notGate[680] ) /* synthesis syn_module_defined=1 */ ;
    input \notGate[679]_keep ;
    output \notGate[680] ;
    
    wire \notGate[679]_keep  /* synthesis alspreserve=1 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(25[15:22])
    
    LUT4 I1 (.A(\notGate[679]_keep ), .B(\notGate[679]_keep ), .C(\notGate[679]_keep ), 
         .D(\notGate[679]_keep ), .Z(\notGate[680] )) /* synthesis syn_instantiated=1, lut_function=((!D !C !B !A)+(!D !C !B A)+(!D !C B !A)+(!D !C B A)+(!D C !B !A)+(!D C !B A)+(!D C B !A)+(!D C B A)), LSE_LINE_FILE_ID=3, LSE_LCOL=13, LSE_RCOL=44, LSE_LLINE=32, LSE_RLINE=32 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(11[2:53])
    defparam I1.init = 16'b0000000011111111;
    
endmodule
//
// Verilog Description of module inverter_U355
//

module inverter_U355 (\notGate[66]_keep , \notGate[67] ) /* synthesis syn_module_defined=1 */ ;
    input \notGate[66]_keep ;
    output \notGate[67] ;
    
    wire \notGate[66]_keep  /* synthesis alspreserve=1 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(25[15:22])
    
    LUT4 I1 (.A(\notGate[66]_keep ), .B(\notGate[66]_keep ), .C(\notGate[66]_keep ), 
         .D(\notGate[66]_keep ), .Z(\notGate[67] )) /* synthesis syn_instantiated=1, lut_function=((!D !C !B !A)+(!D !C !B A)+(!D !C B !A)+(!D !C B A)+(!D C !B !A)+(!D C !B A)+(!D C B !A)+(!D C B A)), LSE_LINE_FILE_ID=3, LSE_LCOL=13, LSE_RCOL=44, LSE_LLINE=32, LSE_RLINE=32 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(11[2:53])
    defparam I1.init = 16'b0000000011111111;
    
endmodule
//
// Verilog Description of module inverter_U356
//

module inverter_U356 (\notGate[678]_keep , \notGate[679] ) /* synthesis syn_module_defined=1 */ ;
    input \notGate[678]_keep ;
    output \notGate[679] ;
    
    wire \notGate[678]_keep  /* synthesis alspreserve=1 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(25[15:22])
    
    LUT4 I1 (.A(\notGate[678]_keep ), .B(\notGate[678]_keep ), .C(\notGate[678]_keep ), 
         .D(\notGate[678]_keep ), .Z(\notGate[679] )) /* synthesis syn_instantiated=1, lut_function=((!D !C !B !A)+(!D !C !B A)+(!D !C B !A)+(!D !C B A)+(!D C !B !A)+(!D C !B A)+(!D C B !A)+(!D C B A)), LSE_LINE_FILE_ID=3, LSE_LCOL=13, LSE_RCOL=44, LSE_LLINE=32, LSE_RLINE=32 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(11[2:53])
    defparam I1.init = 16'b0000000011111111;
    
endmodule
//
// Verilog Description of module inverter_U357
//

module inverter_U357 (\notGate[677]_keep , \notGate[678] ) /* synthesis syn_module_defined=1 */ ;
    input \notGate[677]_keep ;
    output \notGate[678] ;
    
    wire \notGate[677]_keep  /* synthesis alspreserve=1 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(25[15:22])
    
    LUT4 I1 (.A(\notGate[677]_keep ), .B(\notGate[677]_keep ), .C(\notGate[677]_keep ), 
         .D(\notGate[677]_keep ), .Z(\notGate[678] )) /* synthesis syn_instantiated=1, lut_function=((!D !C !B !A)+(!D !C !B A)+(!D !C B !A)+(!D !C B A)+(!D C !B !A)+(!D C !B A)+(!D C B !A)+(!D C B A)), LSE_LINE_FILE_ID=3, LSE_LCOL=13, LSE_RCOL=44, LSE_LLINE=32, LSE_RLINE=32 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(11[2:53])
    defparam I1.init = 16'b0000000011111111;
    
endmodule
//
// Verilog Description of module inverter_U358
//

module inverter_U358 (\notGate[676]_keep , \notGate[677] ) /* synthesis syn_module_defined=1 */ ;
    input \notGate[676]_keep ;
    output \notGate[677] ;
    
    wire \notGate[676]_keep  /* synthesis alspreserve=1 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(25[15:22])
    
    LUT4 I1 (.A(\notGate[676]_keep ), .B(\notGate[676]_keep ), .C(\notGate[676]_keep ), 
         .D(\notGate[676]_keep ), .Z(\notGate[677] )) /* synthesis syn_instantiated=1, lut_function=((!D !C !B !A)+(!D !C !B A)+(!D !C B !A)+(!D !C B A)+(!D C !B !A)+(!D C !B A)+(!D C B !A)+(!D C B A)), LSE_LINE_FILE_ID=3, LSE_LCOL=13, LSE_RCOL=44, LSE_LLINE=32, LSE_RLINE=32 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(11[2:53])
    defparam I1.init = 16'b0000000011111111;
    
endmodule
//
// Verilog Description of module inverter_U359
//

module inverter_U359 (\notGate[675]_keep , \notGate[676] ) /* synthesis syn_module_defined=1 */ ;
    input \notGate[675]_keep ;
    output \notGate[676] ;
    
    wire \notGate[675]_keep  /* synthesis alspreserve=1 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(25[15:22])
    
    LUT4 I1 (.A(\notGate[675]_keep ), .B(\notGate[675]_keep ), .C(\notGate[675]_keep ), 
         .D(\notGate[675]_keep ), .Z(\notGate[676] )) /* synthesis syn_instantiated=1, lut_function=((!D !C !B !A)+(!D !C !B A)+(!D !C B !A)+(!D !C B A)+(!D C !B !A)+(!D C !B A)+(!D C B !A)+(!D C B A)), LSE_LINE_FILE_ID=3, LSE_LCOL=13, LSE_RCOL=44, LSE_LLINE=32, LSE_RLINE=32 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(11[2:53])
    defparam I1.init = 16'b0000000011111111;
    
endmodule
//
// Verilog Description of module inverter_U360
//

module inverter_U360 (\notGate[674]_keep , \notGate[675] ) /* synthesis syn_module_defined=1 */ ;
    input \notGate[674]_keep ;
    output \notGate[675] ;
    
    wire \notGate[674]_keep  /* synthesis alspreserve=1 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(25[15:22])
    
    LUT4 I1 (.A(\notGate[674]_keep ), .B(\notGate[674]_keep ), .C(\notGate[674]_keep ), 
         .D(\notGate[674]_keep ), .Z(\notGate[675] )) /* synthesis syn_instantiated=1, lut_function=((!D !C !B !A)+(!D !C !B A)+(!D !C B !A)+(!D !C B A)+(!D C !B !A)+(!D C !B A)+(!D C B !A)+(!D C B A)), LSE_LINE_FILE_ID=3, LSE_LCOL=13, LSE_RCOL=44, LSE_LLINE=32, LSE_RLINE=32 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(11[2:53])
    defparam I1.init = 16'b0000000011111111;
    
endmodule
//
// Verilog Description of module inverter_U361
//

module inverter_U361 (\notGate[673]_keep , \notGate[674] ) /* synthesis syn_module_defined=1 */ ;
    input \notGate[673]_keep ;
    output \notGate[674] ;
    
    wire \notGate[673]_keep  /* synthesis alspreserve=1 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(25[15:22])
    
    LUT4 I1 (.A(\notGate[673]_keep ), .B(\notGate[673]_keep ), .C(\notGate[673]_keep ), 
         .D(\notGate[673]_keep ), .Z(\notGate[674] )) /* synthesis syn_instantiated=1, lut_function=((!D !C !B !A)+(!D !C !B A)+(!D !C B !A)+(!D !C B A)+(!D C !B !A)+(!D C !B A)+(!D C B !A)+(!D C B A)), LSE_LINE_FILE_ID=3, LSE_LCOL=13, LSE_RCOL=44, LSE_LLINE=32, LSE_RLINE=32 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(11[2:53])
    defparam I1.init = 16'b0000000011111111;
    
endmodule
//
// Verilog Description of module inverter_U362
//

module inverter_U362 (\notGate[672]_keep , \notGate[673] ) /* synthesis syn_module_defined=1 */ ;
    input \notGate[672]_keep ;
    output \notGate[673] ;
    
    wire \notGate[672]_keep  /* synthesis alspreserve=1 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(25[15:22])
    
    LUT4 I1 (.A(\notGate[672]_keep ), .B(\notGate[672]_keep ), .C(\notGate[672]_keep ), 
         .D(\notGate[672]_keep ), .Z(\notGate[673] )) /* synthesis syn_instantiated=1, lut_function=((!D !C !B !A)+(!D !C !B A)+(!D !C B !A)+(!D !C B A)+(!D C !B !A)+(!D C !B A)+(!D C B !A)+(!D C B A)), LSE_LINE_FILE_ID=3, LSE_LCOL=13, LSE_RCOL=44, LSE_LLINE=32, LSE_RLINE=32 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(11[2:53])
    defparam I1.init = 16'b0000000011111111;
    
endmodule
//
// Verilog Description of module inverter_U363
//

module inverter_U363 (\notGate[671]_keep , \notGate[672] ) /* synthesis syn_module_defined=1 */ ;
    input \notGate[671]_keep ;
    output \notGate[672] ;
    
    wire \notGate[671]_keep  /* synthesis alspreserve=1 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(25[15:22])
    
    LUT4 I1 (.A(\notGate[671]_keep ), .B(\notGate[671]_keep ), .C(\notGate[671]_keep ), 
         .D(\notGate[671]_keep ), .Z(\notGate[672] )) /* synthesis syn_instantiated=1, lut_function=((!D !C !B !A)+(!D !C !B A)+(!D !C B !A)+(!D !C B A)+(!D C !B !A)+(!D C !B A)+(!D C B !A)+(!D C B A)), LSE_LINE_FILE_ID=3, LSE_LCOL=13, LSE_RCOL=44, LSE_LLINE=32, LSE_RLINE=32 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(11[2:53])
    defparam I1.init = 16'b0000000011111111;
    
endmodule
//
// Verilog Description of module inverter_U364
//

module inverter_U364 (\notGate[670]_keep , \notGate[671] ) /* synthesis syn_module_defined=1 */ ;
    input \notGate[670]_keep ;
    output \notGate[671] ;
    
    wire \notGate[670]_keep  /* synthesis alspreserve=1 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(25[15:22])
    
    LUT4 I1 (.A(\notGate[670]_keep ), .B(\notGate[670]_keep ), .C(\notGate[670]_keep ), 
         .D(\notGate[670]_keep ), .Z(\notGate[671] )) /* synthesis syn_instantiated=1, lut_function=((!D !C !B !A)+(!D !C !B A)+(!D !C B !A)+(!D !C B A)+(!D C !B !A)+(!D C !B A)+(!D C B !A)+(!D C B A)), LSE_LINE_FILE_ID=3, LSE_LCOL=13, LSE_RCOL=44, LSE_LLINE=32, LSE_RLINE=32 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(11[2:53])
    defparam I1.init = 16'b0000000011111111;
    
endmodule
//
// Verilog Description of module inverter_U365
//

module inverter_U365 (\notGate[669]_keep , \notGate[670] ) /* synthesis syn_module_defined=1 */ ;
    input \notGate[669]_keep ;
    output \notGate[670] ;
    
    wire \notGate[669]_keep  /* synthesis alspreserve=1 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(25[15:22])
    
    LUT4 I1 (.A(\notGate[669]_keep ), .B(\notGate[669]_keep ), .C(\notGate[669]_keep ), 
         .D(\notGate[669]_keep ), .Z(\notGate[670] )) /* synthesis syn_instantiated=1, lut_function=((!D !C !B !A)+(!D !C !B A)+(!D !C B !A)+(!D !C B A)+(!D C !B !A)+(!D C !B A)+(!D C B !A)+(!D C B A)), LSE_LINE_FILE_ID=3, LSE_LCOL=13, LSE_RCOL=44, LSE_LLINE=32, LSE_RLINE=32 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(11[2:53])
    defparam I1.init = 16'b0000000011111111;
    
endmodule
//
// Verilog Description of module inverter_U366
//

module inverter_U366 (\notGate[65]_keep , \notGate[66] ) /* synthesis syn_module_defined=1 */ ;
    input \notGate[65]_keep ;
    output \notGate[66] ;
    
    wire \notGate[65]_keep  /* synthesis alspreserve=1 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(25[15:22])
    
    LUT4 I1 (.A(\notGate[65]_keep ), .B(\notGate[65]_keep ), .C(\notGate[65]_keep ), 
         .D(\notGate[65]_keep ), .Z(\notGate[66] )) /* synthesis syn_instantiated=1, lut_function=((!D !C !B !A)+(!D !C !B A)+(!D !C B !A)+(!D !C B A)+(!D C !B !A)+(!D C !B A)+(!D C B !A)+(!D C B A)), LSE_LINE_FILE_ID=3, LSE_LCOL=13, LSE_RCOL=44, LSE_LLINE=32, LSE_RLINE=32 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(11[2:53])
    defparam I1.init = 16'b0000000011111111;
    
endmodule
//
// Verilog Description of module inverter_U367
//

module inverter_U367 (\notGate[668]_keep , \notGate[669] ) /* synthesis syn_module_defined=1 */ ;
    input \notGate[668]_keep ;
    output \notGate[669] ;
    
    wire \notGate[668]_keep  /* synthesis alspreserve=1 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(25[15:22])
    
    LUT4 I1 (.A(\notGate[668]_keep ), .B(\notGate[668]_keep ), .C(\notGate[668]_keep ), 
         .D(\notGate[668]_keep ), .Z(\notGate[669] )) /* synthesis syn_instantiated=1, lut_function=((!D !C !B !A)+(!D !C !B A)+(!D !C B !A)+(!D !C B A)+(!D C !B !A)+(!D C !B A)+(!D C B !A)+(!D C B A)), LSE_LINE_FILE_ID=3, LSE_LCOL=13, LSE_RCOL=44, LSE_LLINE=32, LSE_RLINE=32 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(11[2:53])
    defparam I1.init = 16'b0000000011111111;
    
endmodule
//
// Verilog Description of module inverter_U368
//

module inverter_U368 (\notGate[667]_keep , \notGate[668] ) /* synthesis syn_module_defined=1 */ ;
    input \notGate[667]_keep ;
    output \notGate[668] ;
    
    wire \notGate[667]_keep  /* synthesis alspreserve=1 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(25[15:22])
    
    LUT4 I1 (.A(\notGate[667]_keep ), .B(\notGate[667]_keep ), .C(\notGate[667]_keep ), 
         .D(\notGate[667]_keep ), .Z(\notGate[668] )) /* synthesis syn_instantiated=1, lut_function=((!D !C !B !A)+(!D !C !B A)+(!D !C B !A)+(!D !C B A)+(!D C !B !A)+(!D C !B A)+(!D C B !A)+(!D C B A)), LSE_LINE_FILE_ID=3, LSE_LCOL=13, LSE_RCOL=44, LSE_LLINE=32, LSE_RLINE=32 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(11[2:53])
    defparam I1.init = 16'b0000000011111111;
    
endmodule
//
// Verilog Description of module inverter_U369
//

module inverter_U369 (\notGate[666]_keep , \notGate[667] ) /* synthesis syn_module_defined=1 */ ;
    input \notGate[666]_keep ;
    output \notGate[667] ;
    
    wire \notGate[666]_keep  /* synthesis alspreserve=1 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(25[15:22])
    
    LUT4 I1 (.A(\notGate[666]_keep ), .B(\notGate[666]_keep ), .C(\notGate[666]_keep ), 
         .D(\notGate[666]_keep ), .Z(\notGate[667] )) /* synthesis syn_instantiated=1, lut_function=((!D !C !B !A)+(!D !C !B A)+(!D !C B !A)+(!D !C B A)+(!D C !B !A)+(!D C !B A)+(!D C B !A)+(!D C B A)), LSE_LINE_FILE_ID=3, LSE_LCOL=13, LSE_RCOL=44, LSE_LLINE=32, LSE_RLINE=32 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(11[2:53])
    defparam I1.init = 16'b0000000011111111;
    
endmodule
//
// Verilog Description of module inverter_U370
//

module inverter_U370 (\notGate[665]_keep , \notGate[666] ) /* synthesis syn_module_defined=1 */ ;
    input \notGate[665]_keep ;
    output \notGate[666] ;
    
    wire \notGate[665]_keep  /* synthesis alspreserve=1 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(25[15:22])
    
    LUT4 I1 (.A(\notGate[665]_keep ), .B(\notGate[665]_keep ), .C(\notGate[665]_keep ), 
         .D(\notGate[665]_keep ), .Z(\notGate[666] )) /* synthesis syn_instantiated=1, lut_function=((!D !C !B !A)+(!D !C !B A)+(!D !C B !A)+(!D !C B A)+(!D C !B !A)+(!D C !B A)+(!D C B !A)+(!D C B A)), LSE_LINE_FILE_ID=3, LSE_LCOL=13, LSE_RCOL=44, LSE_LLINE=32, LSE_RLINE=32 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(11[2:53])
    defparam I1.init = 16'b0000000011111111;
    
endmodule
//
// Verilog Description of module inverter_U371
//

module inverter_U371 (\notGate[664]_keep , \notGate[665] ) /* synthesis syn_module_defined=1 */ ;
    input \notGate[664]_keep ;
    output \notGate[665] ;
    
    wire \notGate[664]_keep  /* synthesis alspreserve=1 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(25[15:22])
    
    LUT4 I1 (.A(\notGate[664]_keep ), .B(\notGate[664]_keep ), .C(\notGate[664]_keep ), 
         .D(\notGate[664]_keep ), .Z(\notGate[665] )) /* synthesis syn_instantiated=1, lut_function=((!D !C !B !A)+(!D !C !B A)+(!D !C B !A)+(!D !C B A)+(!D C !B !A)+(!D C !B A)+(!D C B !A)+(!D C B A)), LSE_LINE_FILE_ID=3, LSE_LCOL=13, LSE_RCOL=44, LSE_LLINE=32, LSE_RLINE=32 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(11[2:53])
    defparam I1.init = 16'b0000000011111111;
    
endmodule
//
// Verilog Description of module inverter_U372
//

module inverter_U372 (\notGate[663]_keep , \notGate[664] ) /* synthesis syn_module_defined=1 */ ;
    input \notGate[663]_keep ;
    output \notGate[664] ;
    
    wire \notGate[663]_keep  /* synthesis alspreserve=1 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(25[15:22])
    
    LUT4 I1 (.A(\notGate[663]_keep ), .B(\notGate[663]_keep ), .C(\notGate[663]_keep ), 
         .D(\notGate[663]_keep ), .Z(\notGate[664] )) /* synthesis syn_instantiated=1, lut_function=((!D !C !B !A)+(!D !C !B A)+(!D !C B !A)+(!D !C B A)+(!D C !B !A)+(!D C !B A)+(!D C B !A)+(!D C B A)), LSE_LINE_FILE_ID=3, LSE_LCOL=13, LSE_RCOL=44, LSE_LLINE=32, LSE_RLINE=32 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(11[2:53])
    defparam I1.init = 16'b0000000011111111;
    
endmodule
//
// Verilog Description of module inverter_U373
//

module inverter_U373 (\notGate[662]_keep , \notGate[663] ) /* synthesis syn_module_defined=1 */ ;
    input \notGate[662]_keep ;
    output \notGate[663] ;
    
    wire \notGate[662]_keep  /* synthesis alspreserve=1 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(25[15:22])
    
    LUT4 I1 (.A(\notGate[662]_keep ), .B(\notGate[662]_keep ), .C(\notGate[662]_keep ), 
         .D(\notGate[662]_keep ), .Z(\notGate[663] )) /* synthesis syn_instantiated=1, lut_function=((!D !C !B !A)+(!D !C !B A)+(!D !C B !A)+(!D !C B A)+(!D C !B !A)+(!D C !B A)+(!D C B !A)+(!D C B A)), LSE_LINE_FILE_ID=3, LSE_LCOL=13, LSE_RCOL=44, LSE_LLINE=32, LSE_RLINE=32 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(11[2:53])
    defparam I1.init = 16'b0000000011111111;
    
endmodule
//
// Verilog Description of module inverter_U374
//

module inverter_U374 (\notGate[661]_keep , \notGate[662] ) /* synthesis syn_module_defined=1 */ ;
    input \notGate[661]_keep ;
    output \notGate[662] ;
    
    wire \notGate[661]_keep  /* synthesis alspreserve=1 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(25[15:22])
    
    LUT4 I1 (.A(\notGate[661]_keep ), .B(\notGate[661]_keep ), .C(\notGate[661]_keep ), 
         .D(\notGate[661]_keep ), .Z(\notGate[662] )) /* synthesis syn_instantiated=1, lut_function=((!D !C !B !A)+(!D !C !B A)+(!D !C B !A)+(!D !C B A)+(!D C !B !A)+(!D C !B A)+(!D C B !A)+(!D C B A)), LSE_LINE_FILE_ID=3, LSE_LCOL=13, LSE_RCOL=44, LSE_LLINE=32, LSE_RLINE=32 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(11[2:53])
    defparam I1.init = 16'b0000000011111111;
    
endmodule
//
// Verilog Description of module inverter_U375
//

module inverter_U375 (\notGate[660]_keep , \notGate[661] ) /* synthesis syn_module_defined=1 */ ;
    input \notGate[660]_keep ;
    output \notGate[661] ;
    
    wire \notGate[660]_keep  /* synthesis alspreserve=1 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(25[15:22])
    
    LUT4 I1 (.A(\notGate[660]_keep ), .B(\notGate[660]_keep ), .C(\notGate[660]_keep ), 
         .D(\notGate[660]_keep ), .Z(\notGate[661] )) /* synthesis syn_instantiated=1, lut_function=((!D !C !B !A)+(!D !C !B A)+(!D !C B !A)+(!D !C B A)+(!D C !B !A)+(!D C !B A)+(!D C B !A)+(!D C B A)), LSE_LINE_FILE_ID=3, LSE_LCOL=13, LSE_RCOL=44, LSE_LLINE=32, LSE_RLINE=32 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(11[2:53])
    defparam I1.init = 16'b0000000011111111;
    
endmodule
//
// Verilog Description of module inverter_U376
//

module inverter_U376 (\notGate[659]_keep , \notGate[660] ) /* synthesis syn_module_defined=1 */ ;
    input \notGate[659]_keep ;
    output \notGate[660] ;
    
    wire \notGate[659]_keep  /* synthesis alspreserve=1 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(25[15:22])
    
    LUT4 I1 (.A(\notGate[659]_keep ), .B(\notGate[659]_keep ), .C(\notGate[659]_keep ), 
         .D(\notGate[659]_keep ), .Z(\notGate[660] )) /* synthesis syn_instantiated=1, lut_function=((!D !C !B !A)+(!D !C !B A)+(!D !C B !A)+(!D !C B A)+(!D C !B !A)+(!D C !B A)+(!D C B !A)+(!D C B A)), LSE_LINE_FILE_ID=3, LSE_LCOL=13, LSE_RCOL=44, LSE_LLINE=32, LSE_RLINE=32 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(11[2:53])
    defparam I1.init = 16'b0000000011111111;
    
endmodule
//
// Verilog Description of module inverter_U377
//

module inverter_U377 (\notGate[64]_keep , \notGate[65] ) /* synthesis syn_module_defined=1 */ ;
    input \notGate[64]_keep ;
    output \notGate[65] ;
    
    wire \notGate[64]_keep  /* synthesis alspreserve=1 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(25[15:22])
    
    LUT4 I1 (.A(\notGate[64]_keep ), .B(\notGate[64]_keep ), .C(\notGate[64]_keep ), 
         .D(\notGate[64]_keep ), .Z(\notGate[65] )) /* synthesis syn_instantiated=1, lut_function=((!D !C !B !A)+(!D !C !B A)+(!D !C B !A)+(!D !C B A)+(!D C !B !A)+(!D C !B A)+(!D C B !A)+(!D C B A)), LSE_LINE_FILE_ID=3, LSE_LCOL=13, LSE_RCOL=44, LSE_LLINE=32, LSE_RLINE=32 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(11[2:53])
    defparam I1.init = 16'b0000000011111111;
    
endmodule
//
// Verilog Description of module inverter_U378
//

module inverter_U378 (\notGate[658]_keep , \notGate[659] ) /* synthesis syn_module_defined=1 */ ;
    input \notGate[658]_keep ;
    output \notGate[659] ;
    
    wire \notGate[658]_keep  /* synthesis alspreserve=1 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(25[15:22])
    
    LUT4 I1 (.A(\notGate[658]_keep ), .B(\notGate[658]_keep ), .C(\notGate[658]_keep ), 
         .D(\notGate[658]_keep ), .Z(\notGate[659] )) /* synthesis syn_instantiated=1, lut_function=((!D !C !B !A)+(!D !C !B A)+(!D !C B !A)+(!D !C B A)+(!D C !B !A)+(!D C !B A)+(!D C B !A)+(!D C B A)), LSE_LINE_FILE_ID=3, LSE_LCOL=13, LSE_RCOL=44, LSE_LLINE=32, LSE_RLINE=32 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(11[2:53])
    defparam I1.init = 16'b0000000011111111;
    
endmodule
//
// Verilog Description of module inverter_U379
//

module inverter_U379 (\notGate[657]_keep , \notGate[658] ) /* synthesis syn_module_defined=1 */ ;
    input \notGate[657]_keep ;
    output \notGate[658] ;
    
    wire \notGate[657]_keep  /* synthesis alspreserve=1 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(25[15:22])
    
    LUT4 I1 (.A(\notGate[657]_keep ), .B(\notGate[657]_keep ), .C(\notGate[657]_keep ), 
         .D(\notGate[657]_keep ), .Z(\notGate[658] )) /* synthesis syn_instantiated=1, lut_function=((!D !C !B !A)+(!D !C !B A)+(!D !C B !A)+(!D !C B A)+(!D C !B !A)+(!D C !B A)+(!D C B !A)+(!D C B A)), LSE_LINE_FILE_ID=3, LSE_LCOL=13, LSE_RCOL=44, LSE_LLINE=32, LSE_RLINE=32 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(11[2:53])
    defparam I1.init = 16'b0000000011111111;
    
endmodule
//
// Verilog Description of module inverter_U380
//

module inverter_U380 (\notGate[656]_keep , \notGate[657] ) /* synthesis syn_module_defined=1 */ ;
    input \notGate[656]_keep ;
    output \notGate[657] ;
    
    wire \notGate[656]_keep  /* synthesis alspreserve=1 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(25[15:22])
    
    LUT4 I1 (.A(\notGate[656]_keep ), .B(\notGate[656]_keep ), .C(\notGate[656]_keep ), 
         .D(\notGate[656]_keep ), .Z(\notGate[657] )) /* synthesis syn_instantiated=1, lut_function=((!D !C !B !A)+(!D !C !B A)+(!D !C B !A)+(!D !C B A)+(!D C !B !A)+(!D C !B A)+(!D C B !A)+(!D C B A)), LSE_LINE_FILE_ID=3, LSE_LCOL=13, LSE_RCOL=44, LSE_LLINE=32, LSE_RLINE=32 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(11[2:53])
    defparam I1.init = 16'b0000000011111111;
    
endmodule
//
// Verilog Description of module inverter_U381
//

module inverter_U381 (\notGate[655]_keep , \notGate[656] ) /* synthesis syn_module_defined=1 */ ;
    input \notGate[655]_keep ;
    output \notGate[656] ;
    
    wire \notGate[655]_keep  /* synthesis alspreserve=1 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(25[15:22])
    
    LUT4 I1 (.A(\notGate[655]_keep ), .B(\notGate[655]_keep ), .C(\notGate[655]_keep ), 
         .D(\notGate[655]_keep ), .Z(\notGate[656] )) /* synthesis syn_instantiated=1, lut_function=((!D !C !B !A)+(!D !C !B A)+(!D !C B !A)+(!D !C B A)+(!D C !B !A)+(!D C !B A)+(!D C B !A)+(!D C B A)), LSE_LINE_FILE_ID=3, LSE_LCOL=13, LSE_RCOL=44, LSE_LLINE=32, LSE_RLINE=32 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(11[2:53])
    defparam I1.init = 16'b0000000011111111;
    
endmodule
//
// Verilog Description of module inverter_U382
//

module inverter_U382 (\notGate[654]_keep , \notGate[655] ) /* synthesis syn_module_defined=1 */ ;
    input \notGate[654]_keep ;
    output \notGate[655] ;
    
    wire \notGate[654]_keep  /* synthesis alspreserve=1 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(25[15:22])
    
    LUT4 I1 (.A(\notGate[654]_keep ), .B(\notGate[654]_keep ), .C(\notGate[654]_keep ), 
         .D(\notGate[654]_keep ), .Z(\notGate[655] )) /* synthesis syn_instantiated=1, lut_function=((!D !C !B !A)+(!D !C !B A)+(!D !C B !A)+(!D !C B A)+(!D C !B !A)+(!D C !B A)+(!D C B !A)+(!D C B A)), LSE_LINE_FILE_ID=3, LSE_LCOL=13, LSE_RCOL=44, LSE_LLINE=32, LSE_RLINE=32 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(11[2:53])
    defparam I1.init = 16'b0000000011111111;
    
endmodule
//
// Verilog Description of module inverter_U383
//

module inverter_U383 (\notGate[653]_keep , \notGate[654] ) /* synthesis syn_module_defined=1 */ ;
    input \notGate[653]_keep ;
    output \notGate[654] ;
    
    wire \notGate[653]_keep  /* synthesis alspreserve=1 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(25[15:22])
    
    LUT4 I1 (.A(\notGate[653]_keep ), .B(\notGate[653]_keep ), .C(\notGate[653]_keep ), 
         .D(\notGate[653]_keep ), .Z(\notGate[654] )) /* synthesis syn_instantiated=1, lut_function=((!D !C !B !A)+(!D !C !B A)+(!D !C B !A)+(!D !C B A)+(!D C !B !A)+(!D C !B A)+(!D C B !A)+(!D C B A)), LSE_LINE_FILE_ID=3, LSE_LCOL=13, LSE_RCOL=44, LSE_LLINE=32, LSE_RLINE=32 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(11[2:53])
    defparam I1.init = 16'b0000000011111111;
    
endmodule
//
// Verilog Description of module inverter_U384
//

module inverter_U384 (\notGate[652]_keep , \notGate[653] ) /* synthesis syn_module_defined=1 */ ;
    input \notGate[652]_keep ;
    output \notGate[653] ;
    
    wire \notGate[652]_keep  /* synthesis alspreserve=1 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(25[15:22])
    
    LUT4 I1 (.A(\notGate[652]_keep ), .B(\notGate[652]_keep ), .C(\notGate[652]_keep ), 
         .D(\notGate[652]_keep ), .Z(\notGate[653] )) /* synthesis syn_instantiated=1, lut_function=((!D !C !B !A)+(!D !C !B A)+(!D !C B !A)+(!D !C B A)+(!D C !B !A)+(!D C !B A)+(!D C B !A)+(!D C B A)), LSE_LINE_FILE_ID=3, LSE_LCOL=13, LSE_RCOL=44, LSE_LLINE=32, LSE_RLINE=32 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(11[2:53])
    defparam I1.init = 16'b0000000011111111;
    
endmodule
//
// Verilog Description of module inverter_U385
//

module inverter_U385 (\notGate[651]_keep , \notGate[652] ) /* synthesis syn_module_defined=1 */ ;
    input \notGate[651]_keep ;
    output \notGate[652] ;
    
    wire \notGate[651]_keep  /* synthesis alspreserve=1 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(25[15:22])
    
    LUT4 I1 (.A(\notGate[651]_keep ), .B(\notGate[651]_keep ), .C(\notGate[651]_keep ), 
         .D(\notGate[651]_keep ), .Z(\notGate[652] )) /* synthesis syn_instantiated=1, lut_function=((!D !C !B !A)+(!D !C !B A)+(!D !C B !A)+(!D !C B A)+(!D C !B !A)+(!D C !B A)+(!D C B !A)+(!D C B A)), LSE_LINE_FILE_ID=3, LSE_LCOL=13, LSE_RCOL=44, LSE_LLINE=32, LSE_RLINE=32 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(11[2:53])
    defparam I1.init = 16'b0000000011111111;
    
endmodule
//
// Verilog Description of module inverter_U386
//

module inverter_U386 (\notGate[650]_keep , \notGate[651] ) /* synthesis syn_module_defined=1 */ ;
    input \notGate[650]_keep ;
    output \notGate[651] ;
    
    wire \notGate[650]_keep  /* synthesis alspreserve=1 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(25[15:22])
    
    LUT4 I1 (.A(\notGate[650]_keep ), .B(\notGate[650]_keep ), .C(\notGate[650]_keep ), 
         .D(\notGate[650]_keep ), .Z(\notGate[651] )) /* synthesis syn_instantiated=1, lut_function=((!D !C !B !A)+(!D !C !B A)+(!D !C B !A)+(!D !C B A)+(!D C !B !A)+(!D C !B A)+(!D C B !A)+(!D C B A)), LSE_LINE_FILE_ID=3, LSE_LCOL=13, LSE_RCOL=44, LSE_LLINE=32, LSE_RLINE=32 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(11[2:53])
    defparam I1.init = 16'b0000000011111111;
    
endmodule
//
// Verilog Description of module inverter_U387
//

module inverter_U387 (\notGate[649]_keep , \notGate[650] ) /* synthesis syn_module_defined=1 */ ;
    input \notGate[649]_keep ;
    output \notGate[650] ;
    
    wire \notGate[649]_keep  /* synthesis alspreserve=1 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(25[15:22])
    
    LUT4 I1 (.A(\notGate[649]_keep ), .B(\notGate[649]_keep ), .C(\notGate[649]_keep ), 
         .D(\notGate[649]_keep ), .Z(\notGate[650] )) /* synthesis syn_instantiated=1, lut_function=((!D !C !B !A)+(!D !C !B A)+(!D !C B !A)+(!D !C B A)+(!D C !B !A)+(!D C !B A)+(!D C B !A)+(!D C B A)), LSE_LINE_FILE_ID=3, LSE_LCOL=13, LSE_RCOL=44, LSE_LLINE=32, LSE_RLINE=32 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(11[2:53])
    defparam I1.init = 16'b0000000011111111;
    
endmodule
//
// Verilog Description of module inverter_U388
//

module inverter_U388 (\notGate[63]_keep , \notGate[64] ) /* synthesis syn_module_defined=1 */ ;
    input \notGate[63]_keep ;
    output \notGate[64] ;
    
    wire \notGate[63]_keep  /* synthesis alspreserve=1 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(25[15:22])
    
    LUT4 I1 (.A(\notGate[63]_keep ), .B(\notGate[63]_keep ), .C(\notGate[63]_keep ), 
         .D(\notGate[63]_keep ), .Z(\notGate[64] )) /* synthesis syn_instantiated=1, lut_function=((!D !C !B !A)+(!D !C !B A)+(!D !C B !A)+(!D !C B A)+(!D C !B !A)+(!D C !B A)+(!D C B !A)+(!D C B A)), LSE_LINE_FILE_ID=3, LSE_LCOL=13, LSE_RCOL=44, LSE_LLINE=32, LSE_RLINE=32 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(11[2:53])
    defparam I1.init = 16'b0000000011111111;
    
endmodule
//
// Verilog Description of module inverter_U389
//

module inverter_U389 (\notGate[648]_keep , \notGate[649] ) /* synthesis syn_module_defined=1 */ ;
    input \notGate[648]_keep ;
    output \notGate[649] ;
    
    wire \notGate[648]_keep  /* synthesis alspreserve=1 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(25[15:22])
    
    LUT4 I1 (.A(\notGate[648]_keep ), .B(\notGate[648]_keep ), .C(\notGate[648]_keep ), 
         .D(\notGate[648]_keep ), .Z(\notGate[649] )) /* synthesis syn_instantiated=1, lut_function=((!D !C !B !A)+(!D !C !B A)+(!D !C B !A)+(!D !C B A)+(!D C !B !A)+(!D C !B A)+(!D C B !A)+(!D C B A)), LSE_LINE_FILE_ID=3, LSE_LCOL=13, LSE_RCOL=44, LSE_LLINE=32, LSE_RLINE=32 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(11[2:53])
    defparam I1.init = 16'b0000000011111111;
    
endmodule
//
// Verilog Description of module inverter_U390
//

module inverter_U390 (\notGate[647]_keep , \notGate[648] ) /* synthesis syn_module_defined=1 */ ;
    input \notGate[647]_keep ;
    output \notGate[648] ;
    
    wire \notGate[647]_keep  /* synthesis alspreserve=1 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(25[15:22])
    
    LUT4 I1 (.A(\notGate[647]_keep ), .B(\notGate[647]_keep ), .C(\notGate[647]_keep ), 
         .D(\notGate[647]_keep ), .Z(\notGate[648] )) /* synthesis syn_instantiated=1, lut_function=((!D !C !B !A)+(!D !C !B A)+(!D !C B !A)+(!D !C B A)+(!D C !B !A)+(!D C !B A)+(!D C B !A)+(!D C B A)), LSE_LINE_FILE_ID=3, LSE_LCOL=13, LSE_RCOL=44, LSE_LLINE=32, LSE_RLINE=32 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(11[2:53])
    defparam I1.init = 16'b0000000011111111;
    
endmodule
//
// Verilog Description of module inverter_U391
//

module inverter_U391 (\notGate[646]_keep , \notGate[647] ) /* synthesis syn_module_defined=1 */ ;
    input \notGate[646]_keep ;
    output \notGate[647] ;
    
    wire \notGate[646]_keep  /* synthesis alspreserve=1 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(25[15:22])
    
    LUT4 I1 (.A(\notGate[646]_keep ), .B(\notGate[646]_keep ), .C(\notGate[646]_keep ), 
         .D(\notGate[646]_keep ), .Z(\notGate[647] )) /* synthesis syn_instantiated=1, lut_function=((!D !C !B !A)+(!D !C !B A)+(!D !C B !A)+(!D !C B A)+(!D C !B !A)+(!D C !B A)+(!D C B !A)+(!D C B A)), LSE_LINE_FILE_ID=3, LSE_LCOL=13, LSE_RCOL=44, LSE_LLINE=32, LSE_RLINE=32 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(11[2:53])
    defparam I1.init = 16'b0000000011111111;
    
endmodule
//
// Verilog Description of module inverter_U392
//

module inverter_U392 (\notGate[645]_keep , \notGate[646] ) /* synthesis syn_module_defined=1 */ ;
    input \notGate[645]_keep ;
    output \notGate[646] ;
    
    wire \notGate[645]_keep  /* synthesis alspreserve=1 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(25[15:22])
    
    LUT4 I1 (.A(\notGate[645]_keep ), .B(\notGate[645]_keep ), .C(\notGate[645]_keep ), 
         .D(\notGate[645]_keep ), .Z(\notGate[646] )) /* synthesis syn_instantiated=1, lut_function=((!D !C !B !A)+(!D !C !B A)+(!D !C B !A)+(!D !C B A)+(!D C !B !A)+(!D C !B A)+(!D C B !A)+(!D C B A)), LSE_LINE_FILE_ID=3, LSE_LCOL=13, LSE_RCOL=44, LSE_LLINE=32, LSE_RLINE=32 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(11[2:53])
    defparam I1.init = 16'b0000000011111111;
    
endmodule
//
// Verilog Description of module inverter_U393
//

module inverter_U393 (\notGate[644]_keep , \notGate[645] ) /* synthesis syn_module_defined=1 */ ;
    input \notGate[644]_keep ;
    output \notGate[645] ;
    
    wire \notGate[644]_keep  /* synthesis alspreserve=1 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(25[15:22])
    
    LUT4 I1 (.A(\notGate[644]_keep ), .B(\notGate[644]_keep ), .C(\notGate[644]_keep ), 
         .D(\notGate[644]_keep ), .Z(\notGate[645] )) /* synthesis syn_instantiated=1, lut_function=((!D !C !B !A)+(!D !C !B A)+(!D !C B !A)+(!D !C B A)+(!D C !B !A)+(!D C !B A)+(!D C B !A)+(!D C B A)), LSE_LINE_FILE_ID=3, LSE_LCOL=13, LSE_RCOL=44, LSE_LLINE=32, LSE_RLINE=32 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(11[2:53])
    defparam I1.init = 16'b0000000011111111;
    
endmodule
//
// Verilog Description of module inverter_U394
//

module inverter_U394 (\notGate[643]_keep , \notGate[644] ) /* synthesis syn_module_defined=1 */ ;
    input \notGate[643]_keep ;
    output \notGate[644] ;
    
    wire \notGate[643]_keep  /* synthesis alspreserve=1 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(25[15:22])
    
    LUT4 I1 (.A(\notGate[643]_keep ), .B(\notGate[643]_keep ), .C(\notGate[643]_keep ), 
         .D(\notGate[643]_keep ), .Z(\notGate[644] )) /* synthesis syn_instantiated=1, lut_function=((!D !C !B !A)+(!D !C !B A)+(!D !C B !A)+(!D !C B A)+(!D C !B !A)+(!D C !B A)+(!D C B !A)+(!D C B A)), LSE_LINE_FILE_ID=3, LSE_LCOL=13, LSE_RCOL=44, LSE_LLINE=32, LSE_RLINE=32 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(11[2:53])
    defparam I1.init = 16'b0000000011111111;
    
endmodule
//
// Verilog Description of module inverter_U395
//

module inverter_U395 (\notGate[642]_keep , \notGate[643] ) /* synthesis syn_module_defined=1 */ ;
    input \notGate[642]_keep ;
    output \notGate[643] ;
    
    wire \notGate[642]_keep  /* synthesis alspreserve=1 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(25[15:22])
    
    LUT4 I1 (.A(\notGate[642]_keep ), .B(\notGate[642]_keep ), .C(\notGate[642]_keep ), 
         .D(\notGate[642]_keep ), .Z(\notGate[643] )) /* synthesis syn_instantiated=1, lut_function=((!D !C !B !A)+(!D !C !B A)+(!D !C B !A)+(!D !C B A)+(!D C !B !A)+(!D C !B A)+(!D C B !A)+(!D C B A)), LSE_LINE_FILE_ID=3, LSE_LCOL=13, LSE_RCOL=44, LSE_LLINE=32, LSE_RLINE=32 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(11[2:53])
    defparam I1.init = 16'b0000000011111111;
    
endmodule
//
// Verilog Description of module inverter_U396
//

module inverter_U396 (\notGate[641]_keep , \notGate[642] ) /* synthesis syn_module_defined=1 */ ;
    input \notGate[641]_keep ;
    output \notGate[642] ;
    
    wire \notGate[641]_keep  /* synthesis alspreserve=1 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(25[15:22])
    
    LUT4 I1 (.A(\notGate[641]_keep ), .B(\notGate[641]_keep ), .C(\notGate[641]_keep ), 
         .D(\notGate[641]_keep ), .Z(\notGate[642] )) /* synthesis syn_instantiated=1, lut_function=((!D !C !B !A)+(!D !C !B A)+(!D !C B !A)+(!D !C B A)+(!D C !B !A)+(!D C !B A)+(!D C B !A)+(!D C B A)), LSE_LINE_FILE_ID=3, LSE_LCOL=13, LSE_RCOL=44, LSE_LLINE=32, LSE_RLINE=32 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(11[2:53])
    defparam I1.init = 16'b0000000011111111;
    
endmodule
//
// Verilog Description of module inverter_U397
//

module inverter_U397 (\notGate[640]_keep , \notGate[641] ) /* synthesis syn_module_defined=1 */ ;
    input \notGate[640]_keep ;
    output \notGate[641] ;
    
    wire \notGate[640]_keep  /* synthesis alspreserve=1 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(25[15:22])
    
    LUT4 I1 (.A(\notGate[640]_keep ), .B(\notGate[640]_keep ), .C(\notGate[640]_keep ), 
         .D(\notGate[640]_keep ), .Z(\notGate[641] )) /* synthesis syn_instantiated=1, lut_function=((!D !C !B !A)+(!D !C !B A)+(!D !C B !A)+(!D !C B A)+(!D C !B !A)+(!D C !B A)+(!D C B !A)+(!D C B A)), LSE_LINE_FILE_ID=3, LSE_LCOL=13, LSE_RCOL=44, LSE_LLINE=32, LSE_RLINE=32 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(11[2:53])
    defparam I1.init = 16'b0000000011111111;
    
endmodule
//
// Verilog Description of module inverter_U398
//

module inverter_U398 (\notGate[639]_keep , \notGate[640] ) /* synthesis syn_module_defined=1 */ ;
    input \notGate[639]_keep ;
    output \notGate[640] ;
    
    wire \notGate[639]_keep  /* synthesis alspreserve=1 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(25[15:22])
    
    LUT4 I1 (.A(\notGate[639]_keep ), .B(\notGate[639]_keep ), .C(\notGate[639]_keep ), 
         .D(\notGate[639]_keep ), .Z(\notGate[640] )) /* synthesis syn_instantiated=1, lut_function=((!D !C !B !A)+(!D !C !B A)+(!D !C B !A)+(!D !C B A)+(!D C !B !A)+(!D C !B A)+(!D C B !A)+(!D C B A)), LSE_LINE_FILE_ID=3, LSE_LCOL=13, LSE_RCOL=44, LSE_LLINE=32, LSE_RLINE=32 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(11[2:53])
    defparam I1.init = 16'b0000000011111111;
    
endmodule
//
// Verilog Description of module inverter_U399
//

module inverter_U399 (\notGate[62]_keep , \notGate[63] ) /* synthesis syn_module_defined=1 */ ;
    input \notGate[62]_keep ;
    output \notGate[63] ;
    
    wire \notGate[62]_keep  /* synthesis alspreserve=1 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(25[15:22])
    
    LUT4 I1 (.A(\notGate[62]_keep ), .B(\notGate[62]_keep ), .C(\notGate[62]_keep ), 
         .D(\notGate[62]_keep ), .Z(\notGate[63] )) /* synthesis syn_instantiated=1, lut_function=((!D !C !B !A)+(!D !C !B A)+(!D !C B !A)+(!D !C B A)+(!D C !B !A)+(!D C !B A)+(!D C B !A)+(!D C B A)), LSE_LINE_FILE_ID=3, LSE_LCOL=13, LSE_RCOL=44, LSE_LLINE=32, LSE_RLINE=32 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(11[2:53])
    defparam I1.init = 16'b0000000011111111;
    
endmodule
//
// Verilog Description of module inverter_U400
//

module inverter_U400 (\notGate[638]_keep , \notGate[639] ) /* synthesis syn_module_defined=1 */ ;
    input \notGate[638]_keep ;
    output \notGate[639] ;
    
    wire \notGate[638]_keep  /* synthesis alspreserve=1 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(25[15:22])
    
    LUT4 I1 (.A(\notGate[638]_keep ), .B(\notGate[638]_keep ), .C(\notGate[638]_keep ), 
         .D(\notGate[638]_keep ), .Z(\notGate[639] )) /* synthesis syn_instantiated=1, lut_function=((!D !C !B !A)+(!D !C !B A)+(!D !C B !A)+(!D !C B A)+(!D C !B !A)+(!D C !B A)+(!D C B !A)+(!D C B A)), LSE_LINE_FILE_ID=3, LSE_LCOL=13, LSE_RCOL=44, LSE_LLINE=32, LSE_RLINE=32 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(11[2:53])
    defparam I1.init = 16'b0000000011111111;
    
endmodule
//
// Verilog Description of module inverter_U401
//

module inverter_U401 (\notGate[637]_keep , \notGate[638] ) /* synthesis syn_module_defined=1 */ ;
    input \notGate[637]_keep ;
    output \notGate[638] ;
    
    wire \notGate[637]_keep  /* synthesis alspreserve=1 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(25[15:22])
    
    LUT4 I1 (.A(\notGate[637]_keep ), .B(\notGate[637]_keep ), .C(\notGate[637]_keep ), 
         .D(\notGate[637]_keep ), .Z(\notGate[638] )) /* synthesis syn_instantiated=1, lut_function=((!D !C !B !A)+(!D !C !B A)+(!D !C B !A)+(!D !C B A)+(!D C !B !A)+(!D C !B A)+(!D C B !A)+(!D C B A)), LSE_LINE_FILE_ID=3, LSE_LCOL=13, LSE_RCOL=44, LSE_LLINE=32, LSE_RLINE=32 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(11[2:53])
    defparam I1.init = 16'b0000000011111111;
    
endmodule
//
// Verilog Description of module inverter_U402
//

module inverter_U402 (\notGate[636]_keep , \notGate[637] ) /* synthesis syn_module_defined=1 */ ;
    input \notGate[636]_keep ;
    output \notGate[637] ;
    
    wire \notGate[636]_keep  /* synthesis alspreserve=1 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(25[15:22])
    
    LUT4 I1 (.A(\notGate[636]_keep ), .B(\notGate[636]_keep ), .C(\notGate[636]_keep ), 
         .D(\notGate[636]_keep ), .Z(\notGate[637] )) /* synthesis syn_instantiated=1, lut_function=((!D !C !B !A)+(!D !C !B A)+(!D !C B !A)+(!D !C B A)+(!D C !B !A)+(!D C !B A)+(!D C B !A)+(!D C B A)), LSE_LINE_FILE_ID=3, LSE_LCOL=13, LSE_RCOL=44, LSE_LLINE=32, LSE_RLINE=32 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(11[2:53])
    defparam I1.init = 16'b0000000011111111;
    
endmodule
//
// Verilog Description of module inverter_U403
//

module inverter_U403 (\notGate[635]_keep , \notGate[636] ) /* synthesis syn_module_defined=1 */ ;
    input \notGate[635]_keep ;
    output \notGate[636] ;
    
    wire \notGate[635]_keep  /* synthesis alspreserve=1 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(25[15:22])
    
    LUT4 I1 (.A(\notGate[635]_keep ), .B(\notGate[635]_keep ), .C(\notGate[635]_keep ), 
         .D(\notGate[635]_keep ), .Z(\notGate[636] )) /* synthesis syn_instantiated=1, lut_function=((!D !C !B !A)+(!D !C !B A)+(!D !C B !A)+(!D !C B A)+(!D C !B !A)+(!D C !B A)+(!D C B !A)+(!D C B A)), LSE_LINE_FILE_ID=3, LSE_LCOL=13, LSE_RCOL=44, LSE_LLINE=32, LSE_RLINE=32 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(11[2:53])
    defparam I1.init = 16'b0000000011111111;
    
endmodule
//
// Verilog Description of module inverter_U404
//

module inverter_U404 (\notGate[634]_keep , \notGate[635] ) /* synthesis syn_module_defined=1 */ ;
    input \notGate[634]_keep ;
    output \notGate[635] ;
    
    wire \notGate[634]_keep  /* synthesis alspreserve=1 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(25[15:22])
    
    LUT4 I1 (.A(\notGate[634]_keep ), .B(\notGate[634]_keep ), .C(\notGate[634]_keep ), 
         .D(\notGate[634]_keep ), .Z(\notGate[635] )) /* synthesis syn_instantiated=1, lut_function=((!D !C !B !A)+(!D !C !B A)+(!D !C B !A)+(!D !C B A)+(!D C !B !A)+(!D C !B A)+(!D C B !A)+(!D C B A)), LSE_LINE_FILE_ID=3, LSE_LCOL=13, LSE_RCOL=44, LSE_LLINE=32, LSE_RLINE=32 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(11[2:53])
    defparam I1.init = 16'b0000000011111111;
    
endmodule
//
// Verilog Description of module inverter_U405
//

module inverter_U405 (\notGate[633]_keep , \notGate[634] ) /* synthesis syn_module_defined=1 */ ;
    input \notGate[633]_keep ;
    output \notGate[634] ;
    
    wire \notGate[633]_keep  /* synthesis alspreserve=1 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(25[15:22])
    
    LUT4 I1 (.A(\notGate[633]_keep ), .B(\notGate[633]_keep ), .C(\notGate[633]_keep ), 
         .D(\notGate[633]_keep ), .Z(\notGate[634] )) /* synthesis syn_instantiated=1, lut_function=((!D !C !B !A)+(!D !C !B A)+(!D !C B !A)+(!D !C B A)+(!D C !B !A)+(!D C !B A)+(!D C B !A)+(!D C B A)), LSE_LINE_FILE_ID=3, LSE_LCOL=13, LSE_RCOL=44, LSE_LLINE=32, LSE_RLINE=32 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(11[2:53])
    defparam I1.init = 16'b0000000011111111;
    
endmodule
//
// Verilog Description of module inverter_U406
//

module inverter_U406 (\notGate[632]_keep , \notGate[633] ) /* synthesis syn_module_defined=1 */ ;
    input \notGate[632]_keep ;
    output \notGate[633] ;
    
    wire \notGate[632]_keep  /* synthesis alspreserve=1 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(25[15:22])
    
    LUT4 I1 (.A(\notGate[632]_keep ), .B(\notGate[632]_keep ), .C(\notGate[632]_keep ), 
         .D(\notGate[632]_keep ), .Z(\notGate[633] )) /* synthesis syn_instantiated=1, lut_function=((!D !C !B !A)+(!D !C !B A)+(!D !C B !A)+(!D !C B A)+(!D C !B !A)+(!D C !B A)+(!D C B !A)+(!D C B A)), LSE_LINE_FILE_ID=3, LSE_LCOL=13, LSE_RCOL=44, LSE_LLINE=32, LSE_RLINE=32 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(11[2:53])
    defparam I1.init = 16'b0000000011111111;
    
endmodule
//
// Verilog Description of module inverter_U407
//

module inverter_U407 (\notGate[631]_keep , \notGate[632] ) /* synthesis syn_module_defined=1 */ ;
    input \notGate[631]_keep ;
    output \notGate[632] ;
    
    wire \notGate[631]_keep  /* synthesis alspreserve=1 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(25[15:22])
    
    LUT4 I1 (.A(\notGate[631]_keep ), .B(\notGate[631]_keep ), .C(\notGate[631]_keep ), 
         .D(\notGate[631]_keep ), .Z(\notGate[632] )) /* synthesis syn_instantiated=1, lut_function=((!D !C !B !A)+(!D !C !B A)+(!D !C B !A)+(!D !C B A)+(!D C !B !A)+(!D C !B A)+(!D C B !A)+(!D C B A)), LSE_LINE_FILE_ID=3, LSE_LCOL=13, LSE_RCOL=44, LSE_LLINE=32, LSE_RLINE=32 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(11[2:53])
    defparam I1.init = 16'b0000000011111111;
    
endmodule
//
// Verilog Description of module inverter_U408
//

module inverter_U408 (\notGate[630]_keep , \notGate[631] ) /* synthesis syn_module_defined=1 */ ;
    input \notGate[630]_keep ;
    output \notGate[631] ;
    
    wire \notGate[630]_keep  /* synthesis alspreserve=1 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(25[15:22])
    
    LUT4 I1 (.A(\notGate[630]_keep ), .B(\notGate[630]_keep ), .C(\notGate[630]_keep ), 
         .D(\notGate[630]_keep ), .Z(\notGate[631] )) /* synthesis syn_instantiated=1, lut_function=((!D !C !B !A)+(!D !C !B A)+(!D !C B !A)+(!D !C B A)+(!D C !B !A)+(!D C !B A)+(!D C B !A)+(!D C B A)), LSE_LINE_FILE_ID=3, LSE_LCOL=13, LSE_RCOL=44, LSE_LLINE=32, LSE_RLINE=32 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(11[2:53])
    defparam I1.init = 16'b0000000011111111;
    
endmodule
//
// Verilog Description of module inverter_U409
//

module inverter_U409 (\notGate[629]_keep , \notGate[630] ) /* synthesis syn_module_defined=1 */ ;
    input \notGate[629]_keep ;
    output \notGate[630] ;
    
    wire \notGate[629]_keep  /* synthesis alspreserve=1 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(25[15:22])
    
    LUT4 I1 (.A(\notGate[629]_keep ), .B(\notGate[629]_keep ), .C(\notGate[629]_keep ), 
         .D(\notGate[629]_keep ), .Z(\notGate[630] )) /* synthesis syn_instantiated=1, lut_function=((!D !C !B !A)+(!D !C !B A)+(!D !C B !A)+(!D !C B A)+(!D C !B !A)+(!D C !B A)+(!D C B !A)+(!D C B A)), LSE_LINE_FILE_ID=3, LSE_LCOL=13, LSE_RCOL=44, LSE_LLINE=32, LSE_RLINE=32 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(11[2:53])
    defparam I1.init = 16'b0000000011111111;
    
endmodule
//
// Verilog Description of module inverter_U410
//

module inverter_U410 (\notGate[61]_keep , \notGate[62] ) /* synthesis syn_module_defined=1 */ ;
    input \notGate[61]_keep ;
    output \notGate[62] ;
    
    wire \notGate[61]_keep  /* synthesis alspreserve=1 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(25[15:22])
    
    LUT4 I1 (.A(\notGate[61]_keep ), .B(\notGate[61]_keep ), .C(\notGate[61]_keep ), 
         .D(\notGate[61]_keep ), .Z(\notGate[62] )) /* synthesis syn_instantiated=1, lut_function=((!D !C !B !A)+(!D !C !B A)+(!D !C B !A)+(!D !C B A)+(!D C !B !A)+(!D C !B A)+(!D C B !A)+(!D C B A)), LSE_LINE_FILE_ID=3, LSE_LCOL=13, LSE_RCOL=44, LSE_LLINE=32, LSE_RLINE=32 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(11[2:53])
    defparam I1.init = 16'b0000000011111111;
    
endmodule
//
// Verilog Description of module inverter_U411
//

module inverter_U411 (\notGate[628]_keep , \notGate[629] ) /* synthesis syn_module_defined=1 */ ;
    input \notGate[628]_keep ;
    output \notGate[629] ;
    
    wire \notGate[628]_keep  /* synthesis alspreserve=1 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(25[15:22])
    
    LUT4 I1 (.A(\notGate[628]_keep ), .B(\notGate[628]_keep ), .C(\notGate[628]_keep ), 
         .D(\notGate[628]_keep ), .Z(\notGate[629] )) /* synthesis syn_instantiated=1, lut_function=((!D !C !B !A)+(!D !C !B A)+(!D !C B !A)+(!D !C B A)+(!D C !B !A)+(!D C !B A)+(!D C B !A)+(!D C B A)), LSE_LINE_FILE_ID=3, LSE_LCOL=13, LSE_RCOL=44, LSE_LLINE=32, LSE_RLINE=32 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(11[2:53])
    defparam I1.init = 16'b0000000011111111;
    
endmodule
//
// Verilog Description of module inverter_U412
//

module inverter_U412 (\notGate[627]_keep , \notGate[628] ) /* synthesis syn_module_defined=1 */ ;
    input \notGate[627]_keep ;
    output \notGate[628] ;
    
    wire \notGate[627]_keep  /* synthesis alspreserve=1 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(25[15:22])
    
    LUT4 I1 (.A(\notGate[627]_keep ), .B(\notGate[627]_keep ), .C(\notGate[627]_keep ), 
         .D(\notGate[627]_keep ), .Z(\notGate[628] )) /* synthesis syn_instantiated=1, lut_function=((!D !C !B !A)+(!D !C !B A)+(!D !C B !A)+(!D !C B A)+(!D C !B !A)+(!D C !B A)+(!D C B !A)+(!D C B A)), LSE_LINE_FILE_ID=3, LSE_LCOL=13, LSE_RCOL=44, LSE_LLINE=32, LSE_RLINE=32 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(11[2:53])
    defparam I1.init = 16'b0000000011111111;
    
endmodule
//
// Verilog Description of module inverter_U413
//

module inverter_U413 (\notGate[626]_keep , \notGate[627] ) /* synthesis syn_module_defined=1 */ ;
    input \notGate[626]_keep ;
    output \notGate[627] ;
    
    wire \notGate[626]_keep  /* synthesis alspreserve=1 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(25[15:22])
    
    LUT4 I1 (.A(\notGate[626]_keep ), .B(\notGate[626]_keep ), .C(\notGate[626]_keep ), 
         .D(\notGate[626]_keep ), .Z(\notGate[627] )) /* synthesis syn_instantiated=1, lut_function=((!D !C !B !A)+(!D !C !B A)+(!D !C B !A)+(!D !C B A)+(!D C !B !A)+(!D C !B A)+(!D C B !A)+(!D C B A)), LSE_LINE_FILE_ID=3, LSE_LCOL=13, LSE_RCOL=44, LSE_LLINE=32, LSE_RLINE=32 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(11[2:53])
    defparam I1.init = 16'b0000000011111111;
    
endmodule
//
// Verilog Description of module inverter_U414
//

module inverter_U414 (\notGate[625]_keep , \notGate[626] ) /* synthesis syn_module_defined=1 */ ;
    input \notGate[625]_keep ;
    output \notGate[626] ;
    
    wire \notGate[625]_keep  /* synthesis alspreserve=1 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(25[15:22])
    
    LUT4 I1 (.A(\notGate[625]_keep ), .B(\notGate[625]_keep ), .C(\notGate[625]_keep ), 
         .D(\notGate[625]_keep ), .Z(\notGate[626] )) /* synthesis syn_instantiated=1, lut_function=((!D !C !B !A)+(!D !C !B A)+(!D !C B !A)+(!D !C B A)+(!D C !B !A)+(!D C !B A)+(!D C B !A)+(!D C B A)), LSE_LINE_FILE_ID=3, LSE_LCOL=13, LSE_RCOL=44, LSE_LLINE=32, LSE_RLINE=32 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(11[2:53])
    defparam I1.init = 16'b0000000011111111;
    
endmodule
//
// Verilog Description of module inverter_U415
//

module inverter_U415 (\notGate[624]_keep , \notGate[625] ) /* synthesis syn_module_defined=1 */ ;
    input \notGate[624]_keep ;
    output \notGate[625] ;
    
    wire \notGate[624]_keep  /* synthesis alspreserve=1 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(25[15:22])
    
    LUT4 I1 (.A(\notGate[624]_keep ), .B(\notGate[624]_keep ), .C(\notGate[624]_keep ), 
         .D(\notGate[624]_keep ), .Z(\notGate[625] )) /* synthesis syn_instantiated=1, lut_function=((!D !C !B !A)+(!D !C !B A)+(!D !C B !A)+(!D !C B A)+(!D C !B !A)+(!D C !B A)+(!D C B !A)+(!D C B A)), LSE_LINE_FILE_ID=3, LSE_LCOL=13, LSE_RCOL=44, LSE_LLINE=32, LSE_RLINE=32 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(11[2:53])
    defparam I1.init = 16'b0000000011111111;
    
endmodule
//
// Verilog Description of module inverter_U416
//

module inverter_U416 (\notGate[623]_keep , \notGate[624] ) /* synthesis syn_module_defined=1 */ ;
    input \notGate[623]_keep ;
    output \notGate[624] ;
    
    wire \notGate[623]_keep  /* synthesis alspreserve=1 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(25[15:22])
    
    LUT4 I1 (.A(\notGate[623]_keep ), .B(\notGate[623]_keep ), .C(\notGate[623]_keep ), 
         .D(\notGate[623]_keep ), .Z(\notGate[624] )) /* synthesis syn_instantiated=1, lut_function=((!D !C !B !A)+(!D !C !B A)+(!D !C B !A)+(!D !C B A)+(!D C !B !A)+(!D C !B A)+(!D C B !A)+(!D C B A)), LSE_LINE_FILE_ID=3, LSE_LCOL=13, LSE_RCOL=44, LSE_LLINE=32, LSE_RLINE=32 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(11[2:53])
    defparam I1.init = 16'b0000000011111111;
    
endmodule
//
// Verilog Description of module inverter_U417
//

module inverter_U417 (\notGate[622]_keep , \notGate[623] ) /* synthesis syn_module_defined=1 */ ;
    input \notGate[622]_keep ;
    output \notGate[623] ;
    
    wire \notGate[622]_keep  /* synthesis alspreserve=1 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(25[15:22])
    
    LUT4 I1 (.A(\notGate[622]_keep ), .B(\notGate[622]_keep ), .C(\notGate[622]_keep ), 
         .D(\notGate[622]_keep ), .Z(\notGate[623] )) /* synthesis syn_instantiated=1, lut_function=((!D !C !B !A)+(!D !C !B A)+(!D !C B !A)+(!D !C B A)+(!D C !B !A)+(!D C !B A)+(!D C B !A)+(!D C B A)), LSE_LINE_FILE_ID=3, LSE_LCOL=13, LSE_RCOL=44, LSE_LLINE=32, LSE_RLINE=32 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(11[2:53])
    defparam I1.init = 16'b0000000011111111;
    
endmodule
//
// Verilog Description of module inverter_U418
//

module inverter_U418 (\notGate[621]_keep , \notGate[622] ) /* synthesis syn_module_defined=1 */ ;
    input \notGate[621]_keep ;
    output \notGate[622] ;
    
    wire \notGate[621]_keep  /* synthesis alspreserve=1 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(25[15:22])
    
    LUT4 I1 (.A(\notGate[621]_keep ), .B(\notGate[621]_keep ), .C(\notGate[621]_keep ), 
         .D(\notGate[621]_keep ), .Z(\notGate[622] )) /* synthesis syn_instantiated=1, lut_function=((!D !C !B !A)+(!D !C !B A)+(!D !C B !A)+(!D !C B A)+(!D C !B !A)+(!D C !B A)+(!D C B !A)+(!D C B A)), LSE_LINE_FILE_ID=3, LSE_LCOL=13, LSE_RCOL=44, LSE_LLINE=32, LSE_RLINE=32 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(11[2:53])
    defparam I1.init = 16'b0000000011111111;
    
endmodule
//
// Verilog Description of module inverter_U419
//

module inverter_U419 (\notGate[620]_keep , \notGate[621] ) /* synthesis syn_module_defined=1 */ ;
    input \notGate[620]_keep ;
    output \notGate[621] ;
    
    wire \notGate[620]_keep  /* synthesis alspreserve=1 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(25[15:22])
    
    LUT4 I1 (.A(\notGate[620]_keep ), .B(\notGate[620]_keep ), .C(\notGate[620]_keep ), 
         .D(\notGate[620]_keep ), .Z(\notGate[621] )) /* synthesis syn_instantiated=1, lut_function=((!D !C !B !A)+(!D !C !B A)+(!D !C B !A)+(!D !C B A)+(!D C !B !A)+(!D C !B A)+(!D C B !A)+(!D C B A)), LSE_LINE_FILE_ID=3, LSE_LCOL=13, LSE_RCOL=44, LSE_LLINE=32, LSE_RLINE=32 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(11[2:53])
    defparam I1.init = 16'b0000000011111111;
    
endmodule
//
// Verilog Description of module inverter_U420
//

module inverter_U420 (\notGate[619]_keep , \notGate[620] ) /* synthesis syn_module_defined=1 */ ;
    input \notGate[619]_keep ;
    output \notGate[620] ;
    
    wire \notGate[619]_keep  /* synthesis alspreserve=1 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(25[15:22])
    
    LUT4 I1 (.A(\notGate[619]_keep ), .B(\notGate[619]_keep ), .C(\notGate[619]_keep ), 
         .D(\notGate[619]_keep ), .Z(\notGate[620] )) /* synthesis syn_instantiated=1, lut_function=((!D !C !B !A)+(!D !C !B A)+(!D !C B !A)+(!D !C B A)+(!D C !B !A)+(!D C !B A)+(!D C B !A)+(!D C B A)), LSE_LINE_FILE_ID=3, LSE_LCOL=13, LSE_RCOL=44, LSE_LLINE=32, LSE_RLINE=32 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(11[2:53])
    defparam I1.init = 16'b0000000011111111;
    
endmodule
//
// Verilog Description of module inverter_U421
//

module inverter_U421 (\notGate[60]_keep , \notGate[61] ) /* synthesis syn_module_defined=1 */ ;
    input \notGate[60]_keep ;
    output \notGate[61] ;
    
    wire \notGate[60]_keep  /* synthesis alspreserve=1 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(25[15:22])
    
    LUT4 I1 (.A(\notGate[60]_keep ), .B(\notGate[60]_keep ), .C(\notGate[60]_keep ), 
         .D(\notGate[60]_keep ), .Z(\notGate[61] )) /* synthesis syn_instantiated=1, lut_function=((!D !C !B !A)+(!D !C !B A)+(!D !C B !A)+(!D !C B A)+(!D C !B !A)+(!D C !B A)+(!D C B !A)+(!D C B A)), LSE_LINE_FILE_ID=3, LSE_LCOL=13, LSE_RCOL=44, LSE_LLINE=32, LSE_RLINE=32 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(11[2:53])
    defparam I1.init = 16'b0000000011111111;
    
endmodule
//
// Verilog Description of module inverter_U422
//

module inverter_U422 (\notGate[618]_keep , \notGate[619] ) /* synthesis syn_module_defined=1 */ ;
    input \notGate[618]_keep ;
    output \notGate[619] ;
    
    wire \notGate[618]_keep  /* synthesis alspreserve=1 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(25[15:22])
    
    LUT4 I1 (.A(\notGate[618]_keep ), .B(\notGate[618]_keep ), .C(\notGate[618]_keep ), 
         .D(\notGate[618]_keep ), .Z(\notGate[619] )) /* synthesis syn_instantiated=1, lut_function=((!D !C !B !A)+(!D !C !B A)+(!D !C B !A)+(!D !C B A)+(!D C !B !A)+(!D C !B A)+(!D C B !A)+(!D C B A)), LSE_LINE_FILE_ID=3, LSE_LCOL=13, LSE_RCOL=44, LSE_LLINE=32, LSE_RLINE=32 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(11[2:53])
    defparam I1.init = 16'b0000000011111111;
    
endmodule
//
// Verilog Description of module inverter_U423
//

module inverter_U423 (\notGate[617]_keep , \notGate[618] ) /* synthesis syn_module_defined=1 */ ;
    input \notGate[617]_keep ;
    output \notGate[618] ;
    
    wire \notGate[617]_keep  /* synthesis alspreserve=1 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(25[15:22])
    
    LUT4 I1 (.A(\notGate[617]_keep ), .B(\notGate[617]_keep ), .C(\notGate[617]_keep ), 
         .D(\notGate[617]_keep ), .Z(\notGate[618] )) /* synthesis syn_instantiated=1, lut_function=((!D !C !B !A)+(!D !C !B A)+(!D !C B !A)+(!D !C B A)+(!D C !B !A)+(!D C !B A)+(!D C B !A)+(!D C B A)), LSE_LINE_FILE_ID=3, LSE_LCOL=13, LSE_RCOL=44, LSE_LLINE=32, LSE_RLINE=32 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(11[2:53])
    defparam I1.init = 16'b0000000011111111;
    
endmodule
//
// Verilog Description of module inverter_U424
//

module inverter_U424 (\notGate[616]_keep , \notGate[617] ) /* synthesis syn_module_defined=1 */ ;
    input \notGate[616]_keep ;
    output \notGate[617] ;
    
    wire \notGate[616]_keep  /* synthesis alspreserve=1 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(25[15:22])
    
    LUT4 I1 (.A(\notGate[616]_keep ), .B(\notGate[616]_keep ), .C(\notGate[616]_keep ), 
         .D(\notGate[616]_keep ), .Z(\notGate[617] )) /* synthesis syn_instantiated=1, lut_function=((!D !C !B !A)+(!D !C !B A)+(!D !C B !A)+(!D !C B A)+(!D C !B !A)+(!D C !B A)+(!D C B !A)+(!D C B A)), LSE_LINE_FILE_ID=3, LSE_LCOL=13, LSE_RCOL=44, LSE_LLINE=32, LSE_RLINE=32 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(11[2:53])
    defparam I1.init = 16'b0000000011111111;
    
endmodule
//
// Verilog Description of module inverter_U425
//

module inverter_U425 (\notGate[615]_keep , \notGate[616] ) /* synthesis syn_module_defined=1 */ ;
    input \notGate[615]_keep ;
    output \notGate[616] ;
    
    wire \notGate[615]_keep  /* synthesis alspreserve=1 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(25[15:22])
    
    LUT4 I1 (.A(\notGate[615]_keep ), .B(\notGate[615]_keep ), .C(\notGate[615]_keep ), 
         .D(\notGate[615]_keep ), .Z(\notGate[616] )) /* synthesis syn_instantiated=1, lut_function=((!D !C !B !A)+(!D !C !B A)+(!D !C B !A)+(!D !C B A)+(!D C !B !A)+(!D C !B A)+(!D C B !A)+(!D C B A)), LSE_LINE_FILE_ID=3, LSE_LCOL=13, LSE_RCOL=44, LSE_LLINE=32, LSE_RLINE=32 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(11[2:53])
    defparam I1.init = 16'b0000000011111111;
    
endmodule
//
// Verilog Description of module inverter_U426
//

module inverter_U426 (\notGate[614]_keep , \notGate[615] ) /* synthesis syn_module_defined=1 */ ;
    input \notGate[614]_keep ;
    output \notGate[615] ;
    
    wire \notGate[614]_keep  /* synthesis alspreserve=1 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(25[15:22])
    
    LUT4 I1 (.A(\notGate[614]_keep ), .B(\notGate[614]_keep ), .C(\notGate[614]_keep ), 
         .D(\notGate[614]_keep ), .Z(\notGate[615] )) /* synthesis syn_instantiated=1, lut_function=((!D !C !B !A)+(!D !C !B A)+(!D !C B !A)+(!D !C B A)+(!D C !B !A)+(!D C !B A)+(!D C B !A)+(!D C B A)), LSE_LINE_FILE_ID=3, LSE_LCOL=13, LSE_RCOL=44, LSE_LLINE=32, LSE_RLINE=32 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(11[2:53])
    defparam I1.init = 16'b0000000011111111;
    
endmodule
//
// Verilog Description of module inverter_U427
//

module inverter_U427 (\notGate[613]_keep , \notGate[614] ) /* synthesis syn_module_defined=1 */ ;
    input \notGate[613]_keep ;
    output \notGate[614] ;
    
    wire \notGate[613]_keep  /* synthesis alspreserve=1 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(25[15:22])
    
    LUT4 I1 (.A(\notGate[613]_keep ), .B(\notGate[613]_keep ), .C(\notGate[613]_keep ), 
         .D(\notGate[613]_keep ), .Z(\notGate[614] )) /* synthesis syn_instantiated=1, lut_function=((!D !C !B !A)+(!D !C !B A)+(!D !C B !A)+(!D !C B A)+(!D C !B !A)+(!D C !B A)+(!D C B !A)+(!D C B A)), LSE_LINE_FILE_ID=3, LSE_LCOL=13, LSE_RCOL=44, LSE_LLINE=32, LSE_RLINE=32 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(11[2:53])
    defparam I1.init = 16'b0000000011111111;
    
endmodule
//
// Verilog Description of module inverter_U428
//

module inverter_U428 (\notGate[612]_keep , \notGate[613] ) /* synthesis syn_module_defined=1 */ ;
    input \notGate[612]_keep ;
    output \notGate[613] ;
    
    wire \notGate[612]_keep  /* synthesis alspreserve=1 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(25[15:22])
    
    LUT4 I1 (.A(\notGate[612]_keep ), .B(\notGate[612]_keep ), .C(\notGate[612]_keep ), 
         .D(\notGate[612]_keep ), .Z(\notGate[613] )) /* synthesis syn_instantiated=1, lut_function=((!D !C !B !A)+(!D !C !B A)+(!D !C B !A)+(!D !C B A)+(!D C !B !A)+(!D C !B A)+(!D C B !A)+(!D C B A)), LSE_LINE_FILE_ID=3, LSE_LCOL=13, LSE_RCOL=44, LSE_LLINE=32, LSE_RLINE=32 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(11[2:53])
    defparam I1.init = 16'b0000000011111111;
    
endmodule
//
// Verilog Description of module inverter_U429
//

module inverter_U429 (\notGate[611]_keep , \notGate[612] ) /* synthesis syn_module_defined=1 */ ;
    input \notGate[611]_keep ;
    output \notGate[612] ;
    
    wire \notGate[611]_keep  /* synthesis alspreserve=1 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(25[15:22])
    
    LUT4 I1 (.A(\notGate[611]_keep ), .B(\notGate[611]_keep ), .C(\notGate[611]_keep ), 
         .D(\notGate[611]_keep ), .Z(\notGate[612] )) /* synthesis syn_instantiated=1, lut_function=((!D !C !B !A)+(!D !C !B A)+(!D !C B !A)+(!D !C B A)+(!D C !B !A)+(!D C !B A)+(!D C B !A)+(!D C B A)), LSE_LINE_FILE_ID=3, LSE_LCOL=13, LSE_RCOL=44, LSE_LLINE=32, LSE_RLINE=32 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(11[2:53])
    defparam I1.init = 16'b0000000011111111;
    
endmodule
//
// Verilog Description of module inverter_U430
//

module inverter_U430 (\notGate[610]_keep , \notGate[611] ) /* synthesis syn_module_defined=1 */ ;
    input \notGate[610]_keep ;
    output \notGate[611] ;
    
    wire \notGate[610]_keep  /* synthesis alspreserve=1 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(25[15:22])
    
    LUT4 I1 (.A(\notGate[610]_keep ), .B(\notGate[610]_keep ), .C(\notGate[610]_keep ), 
         .D(\notGate[610]_keep ), .Z(\notGate[611] )) /* synthesis syn_instantiated=1, lut_function=((!D !C !B !A)+(!D !C !B A)+(!D !C B !A)+(!D !C B A)+(!D C !B !A)+(!D C !B A)+(!D C B !A)+(!D C B A)), LSE_LINE_FILE_ID=3, LSE_LCOL=13, LSE_RCOL=44, LSE_LLINE=32, LSE_RLINE=32 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(11[2:53])
    defparam I1.init = 16'b0000000011111111;
    
endmodule
//
// Verilog Description of module inverter_U431
//

module inverter_U431 (\notGate[609]_keep , \notGate[610] ) /* synthesis syn_module_defined=1 */ ;
    input \notGate[609]_keep ;
    output \notGate[610] ;
    
    wire \notGate[609]_keep  /* synthesis alspreserve=1 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(25[15:22])
    
    LUT4 I1 (.A(\notGate[609]_keep ), .B(\notGate[609]_keep ), .C(\notGate[609]_keep ), 
         .D(\notGate[609]_keep ), .Z(\notGate[610] )) /* synthesis syn_instantiated=1, lut_function=((!D !C !B !A)+(!D !C !B A)+(!D !C B !A)+(!D !C B A)+(!D C !B !A)+(!D C !B A)+(!D C B !A)+(!D C B A)), LSE_LINE_FILE_ID=3, LSE_LCOL=13, LSE_RCOL=44, LSE_LLINE=32, LSE_RLINE=32 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(11[2:53])
    defparam I1.init = 16'b0000000011111111;
    
endmodule
//
// Verilog Description of module inverter_U432
//

module inverter_U432 (\notGate[59]_keep , \notGate[60] ) /* synthesis syn_module_defined=1 */ ;
    input \notGate[59]_keep ;
    output \notGate[60] ;
    
    wire \notGate[59]_keep  /* synthesis alspreserve=1 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(25[15:22])
    
    LUT4 I1 (.A(\notGate[59]_keep ), .B(\notGate[59]_keep ), .C(\notGate[59]_keep ), 
         .D(\notGate[59]_keep ), .Z(\notGate[60] )) /* synthesis syn_instantiated=1, lut_function=((!D !C !B !A)+(!D !C !B A)+(!D !C B !A)+(!D !C B A)+(!D C !B !A)+(!D C !B A)+(!D C B !A)+(!D C B A)), LSE_LINE_FILE_ID=3, LSE_LCOL=13, LSE_RCOL=44, LSE_LLINE=32, LSE_RLINE=32 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(11[2:53])
    defparam I1.init = 16'b0000000011111111;
    
endmodule
//
// Verilog Description of module inverter_U433
//

module inverter_U433 (\notGate[608]_keep , \notGate[609] ) /* synthesis syn_module_defined=1 */ ;
    input \notGate[608]_keep ;
    output \notGate[609] ;
    
    wire \notGate[608]_keep  /* synthesis alspreserve=1 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(25[15:22])
    
    LUT4 I1 (.A(\notGate[608]_keep ), .B(\notGate[608]_keep ), .C(\notGate[608]_keep ), 
         .D(\notGate[608]_keep ), .Z(\notGate[609] )) /* synthesis syn_instantiated=1, lut_function=((!D !C !B !A)+(!D !C !B A)+(!D !C B !A)+(!D !C B A)+(!D C !B !A)+(!D C !B A)+(!D C B !A)+(!D C B A)), LSE_LINE_FILE_ID=3, LSE_LCOL=13, LSE_RCOL=44, LSE_LLINE=32, LSE_RLINE=32 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(11[2:53])
    defparam I1.init = 16'b0000000011111111;
    
endmodule
//
// Verilog Description of module inverter_U434
//

module inverter_U434 (\notGate[607]_keep , \notGate[608] ) /* synthesis syn_module_defined=1 */ ;
    input \notGate[607]_keep ;
    output \notGate[608] ;
    
    wire \notGate[607]_keep  /* synthesis alspreserve=1 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(25[15:22])
    
    LUT4 I1 (.A(\notGate[607]_keep ), .B(\notGate[607]_keep ), .C(\notGate[607]_keep ), 
         .D(\notGate[607]_keep ), .Z(\notGate[608] )) /* synthesis syn_instantiated=1, lut_function=((!D !C !B !A)+(!D !C !B A)+(!D !C B !A)+(!D !C B A)+(!D C !B !A)+(!D C !B A)+(!D C B !A)+(!D C B A)), LSE_LINE_FILE_ID=3, LSE_LCOL=13, LSE_RCOL=44, LSE_LLINE=32, LSE_RLINE=32 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(11[2:53])
    defparam I1.init = 16'b0000000011111111;
    
endmodule
//
// Verilog Description of module inverter_U435
//

module inverter_U435 (\notGate[606]_keep , \notGate[607] ) /* synthesis syn_module_defined=1 */ ;
    input \notGate[606]_keep ;
    output \notGate[607] ;
    
    wire \notGate[606]_keep  /* synthesis alspreserve=1 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(25[15:22])
    
    LUT4 I1 (.A(\notGate[606]_keep ), .B(\notGate[606]_keep ), .C(\notGate[606]_keep ), 
         .D(\notGate[606]_keep ), .Z(\notGate[607] )) /* synthesis syn_instantiated=1, lut_function=((!D !C !B !A)+(!D !C !B A)+(!D !C B !A)+(!D !C B A)+(!D C !B !A)+(!D C !B A)+(!D C B !A)+(!D C B A)), LSE_LINE_FILE_ID=3, LSE_LCOL=13, LSE_RCOL=44, LSE_LLINE=32, LSE_RLINE=32 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(11[2:53])
    defparam I1.init = 16'b0000000011111111;
    
endmodule
//
// Verilog Description of module inverter_U436
//

module inverter_U436 (\notGate[605]_keep , \notGate[606] ) /* synthesis syn_module_defined=1 */ ;
    input \notGate[605]_keep ;
    output \notGate[606] ;
    
    wire \notGate[605]_keep  /* synthesis alspreserve=1 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(25[15:22])
    
    LUT4 I1 (.A(\notGate[605]_keep ), .B(\notGate[605]_keep ), .C(\notGate[605]_keep ), 
         .D(\notGate[605]_keep ), .Z(\notGate[606] )) /* synthesis syn_instantiated=1, lut_function=((!D !C !B !A)+(!D !C !B A)+(!D !C B !A)+(!D !C B A)+(!D C !B !A)+(!D C !B A)+(!D C B !A)+(!D C B A)), LSE_LINE_FILE_ID=3, LSE_LCOL=13, LSE_RCOL=44, LSE_LLINE=32, LSE_RLINE=32 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(11[2:53])
    defparam I1.init = 16'b0000000011111111;
    
endmodule
//
// Verilog Description of module inverter_U437
//

module inverter_U437 (\notGate[604]_keep , \notGate[605] ) /* synthesis syn_module_defined=1 */ ;
    input \notGate[604]_keep ;
    output \notGate[605] ;
    
    wire \notGate[604]_keep  /* synthesis alspreserve=1 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(25[15:22])
    
    LUT4 I1 (.A(\notGate[604]_keep ), .B(\notGate[604]_keep ), .C(\notGate[604]_keep ), 
         .D(\notGate[604]_keep ), .Z(\notGate[605] )) /* synthesis syn_instantiated=1, lut_function=((!D !C !B !A)+(!D !C !B A)+(!D !C B !A)+(!D !C B A)+(!D C !B !A)+(!D C !B A)+(!D C B !A)+(!D C B A)), LSE_LINE_FILE_ID=3, LSE_LCOL=13, LSE_RCOL=44, LSE_LLINE=32, LSE_RLINE=32 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(11[2:53])
    defparam I1.init = 16'b0000000011111111;
    
endmodule
//
// Verilog Description of module inverter_U438
//

module inverter_U438 (\notGate[603]_keep , \notGate[604] ) /* synthesis syn_module_defined=1 */ ;
    input \notGate[603]_keep ;
    output \notGate[604] ;
    
    wire \notGate[603]_keep  /* synthesis alspreserve=1 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(25[15:22])
    
    LUT4 I1 (.A(\notGate[603]_keep ), .B(\notGate[603]_keep ), .C(\notGate[603]_keep ), 
         .D(\notGate[603]_keep ), .Z(\notGate[604] )) /* synthesis syn_instantiated=1, lut_function=((!D !C !B !A)+(!D !C !B A)+(!D !C B !A)+(!D !C B A)+(!D C !B !A)+(!D C !B A)+(!D C B !A)+(!D C B A)), LSE_LINE_FILE_ID=3, LSE_LCOL=13, LSE_RCOL=44, LSE_LLINE=32, LSE_RLINE=32 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(11[2:53])
    defparam I1.init = 16'b0000000011111111;
    
endmodule
//
// Verilog Description of module inverter_U439
//

module inverter_U439 (\notGate[602]_keep , \notGate[603] ) /* synthesis syn_module_defined=1 */ ;
    input \notGate[602]_keep ;
    output \notGate[603] ;
    
    wire \notGate[602]_keep  /* synthesis alspreserve=1 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(25[15:22])
    
    LUT4 I1 (.A(\notGate[602]_keep ), .B(\notGate[602]_keep ), .C(\notGate[602]_keep ), 
         .D(\notGate[602]_keep ), .Z(\notGate[603] )) /* synthesis syn_instantiated=1, lut_function=((!D !C !B !A)+(!D !C !B A)+(!D !C B !A)+(!D !C B A)+(!D C !B !A)+(!D C !B A)+(!D C B !A)+(!D C B A)), LSE_LINE_FILE_ID=3, LSE_LCOL=13, LSE_RCOL=44, LSE_LLINE=32, LSE_RLINE=32 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(11[2:53])
    defparam I1.init = 16'b0000000011111111;
    
endmodule
//
// Verilog Description of module inverter_U440
//

module inverter_U440 (\notGate[601]_keep , \notGate[602] ) /* synthesis syn_module_defined=1 */ ;
    input \notGate[601]_keep ;
    output \notGate[602] ;
    
    wire \notGate[601]_keep  /* synthesis alspreserve=1 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(25[15:22])
    
    LUT4 I1 (.A(\notGate[601]_keep ), .B(\notGate[601]_keep ), .C(\notGate[601]_keep ), 
         .D(\notGate[601]_keep ), .Z(\notGate[602] )) /* synthesis syn_instantiated=1, lut_function=((!D !C !B !A)+(!D !C !B A)+(!D !C B !A)+(!D !C B A)+(!D C !B !A)+(!D C !B A)+(!D C B !A)+(!D C B A)), LSE_LINE_FILE_ID=3, LSE_LCOL=13, LSE_RCOL=44, LSE_LLINE=32, LSE_RLINE=32 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(11[2:53])
    defparam I1.init = 16'b0000000011111111;
    
endmodule
//
// Verilog Description of module inverter_U441
//

module inverter_U441 (\notGate[600]_keep , \notGate[601] ) /* synthesis syn_module_defined=1 */ ;
    input \notGate[600]_keep ;
    output \notGate[601] ;
    
    wire \notGate[600]_keep  /* synthesis alspreserve=1 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(25[15:22])
    
    LUT4 I1 (.A(\notGate[600]_keep ), .B(\notGate[600]_keep ), .C(\notGate[600]_keep ), 
         .D(\notGate[600]_keep ), .Z(\notGate[601] )) /* synthesis syn_instantiated=1, lut_function=((!D !C !B !A)+(!D !C !B A)+(!D !C B !A)+(!D !C B A)+(!D C !B !A)+(!D C !B A)+(!D C B !A)+(!D C B A)), LSE_LINE_FILE_ID=3, LSE_LCOL=13, LSE_RCOL=44, LSE_LLINE=32, LSE_RLINE=32 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(11[2:53])
    defparam I1.init = 16'b0000000011111111;
    
endmodule
//
// Verilog Description of module inverter_U442
//

module inverter_U442 (\notGate[599]_keep , \notGate[600] ) /* synthesis syn_module_defined=1 */ ;
    input \notGate[599]_keep ;
    output \notGate[600] ;
    
    wire \notGate[599]_keep  /* synthesis alspreserve=1 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(25[15:22])
    
    LUT4 I1 (.A(\notGate[599]_keep ), .B(\notGate[599]_keep ), .C(\notGate[599]_keep ), 
         .D(\notGate[599]_keep ), .Z(\notGate[600] )) /* synthesis syn_instantiated=1, lut_function=((!D !C !B !A)+(!D !C !B A)+(!D !C B !A)+(!D !C B A)+(!D C !B !A)+(!D C !B A)+(!D C B !A)+(!D C B A)), LSE_LINE_FILE_ID=3, LSE_LCOL=13, LSE_RCOL=44, LSE_LLINE=32, LSE_RLINE=32 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(11[2:53])
    defparam I1.init = 16'b0000000011111111;
    
endmodule
//
// Verilog Description of module inverter_U443
//

module inverter_U443 (\notGate[4]_keep , \notGate[5] ) /* synthesis syn_module_defined=1 */ ;
    input \notGate[4]_keep ;
    output \notGate[5] ;
    
    wire \notGate[4]_keep  /* synthesis alspreserve=1 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(25[15:22])
    
    LUT4 I1 (.A(\notGate[4]_keep ), .B(\notGate[4]_keep ), .C(\notGate[4]_keep ), 
         .D(\notGate[4]_keep ), .Z(\notGate[5] )) /* synthesis syn_instantiated=1, lut_function=((!D !C !B !A)+(!D !C !B A)+(!D !C B !A)+(!D !C B A)+(!D C !B !A)+(!D C !B A)+(!D C B !A)+(!D C B A)), LSE_LINE_FILE_ID=3, LSE_LCOL=13, LSE_RCOL=44, LSE_LLINE=32, LSE_RLINE=32 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(11[2:53])
    defparam I1.init = 16'b0000000011111111;
    
endmodule
//
// Verilog Description of module inverter_U444
//

module inverter_U444 (\notGate[58]_keep , \notGate[59] ) /* synthesis syn_module_defined=1 */ ;
    input \notGate[58]_keep ;
    output \notGate[59] ;
    
    wire \notGate[58]_keep  /* synthesis alspreserve=1 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(25[15:22])
    
    LUT4 I1 (.A(\notGate[58]_keep ), .B(\notGate[58]_keep ), .C(\notGate[58]_keep ), 
         .D(\notGate[58]_keep ), .Z(\notGate[59] )) /* synthesis syn_instantiated=1, lut_function=((!D !C !B !A)+(!D !C !B A)+(!D !C B !A)+(!D !C B A)+(!D C !B !A)+(!D C !B A)+(!D C B !A)+(!D C B A)), LSE_LINE_FILE_ID=3, LSE_LCOL=13, LSE_RCOL=44, LSE_LLINE=32, LSE_RLINE=32 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(11[2:53])
    defparam I1.init = 16'b0000000011111111;
    
endmodule
//
// Verilog Description of module inverter_U445
//

module inverter_U445 (\notGate[598]_keep , \notGate[599] ) /* synthesis syn_module_defined=1 */ ;
    input \notGate[598]_keep ;
    output \notGate[599] ;
    
    wire \notGate[598]_keep  /* synthesis alspreserve=1 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(25[15:22])
    
    LUT4 I1 (.A(\notGate[598]_keep ), .B(\notGate[598]_keep ), .C(\notGate[598]_keep ), 
         .D(\notGate[598]_keep ), .Z(\notGate[599] )) /* synthesis syn_instantiated=1, lut_function=((!D !C !B !A)+(!D !C !B A)+(!D !C B !A)+(!D !C B A)+(!D C !B !A)+(!D C !B A)+(!D C B !A)+(!D C B A)), LSE_LINE_FILE_ID=3, LSE_LCOL=13, LSE_RCOL=44, LSE_LLINE=32, LSE_RLINE=32 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(11[2:53])
    defparam I1.init = 16'b0000000011111111;
    
endmodule
//
// Verilog Description of module inverter_U446
//

module inverter_U446 (\notGate[597]_keep , \notGate[598] ) /* synthesis syn_module_defined=1 */ ;
    input \notGate[597]_keep ;
    output \notGate[598] ;
    
    wire \notGate[597]_keep  /* synthesis alspreserve=1 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(25[15:22])
    
    LUT4 I1 (.A(\notGate[597]_keep ), .B(\notGate[597]_keep ), .C(\notGate[597]_keep ), 
         .D(\notGate[597]_keep ), .Z(\notGate[598] )) /* synthesis syn_instantiated=1, lut_function=((!D !C !B !A)+(!D !C !B A)+(!D !C B !A)+(!D !C B A)+(!D C !B !A)+(!D C !B A)+(!D C B !A)+(!D C B A)), LSE_LINE_FILE_ID=3, LSE_LCOL=13, LSE_RCOL=44, LSE_LLINE=32, LSE_RLINE=32 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(11[2:53])
    defparam I1.init = 16'b0000000011111111;
    
endmodule
//
// Verilog Description of module inverter_U447
//

module inverter_U447 (\notGate[596]_keep , \notGate[597] ) /* synthesis syn_module_defined=1 */ ;
    input \notGate[596]_keep ;
    output \notGate[597] ;
    
    wire \notGate[596]_keep  /* synthesis alspreserve=1 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(25[15:22])
    
    LUT4 I1 (.A(\notGate[596]_keep ), .B(\notGate[596]_keep ), .C(\notGate[596]_keep ), 
         .D(\notGate[596]_keep ), .Z(\notGate[597] )) /* synthesis syn_instantiated=1, lut_function=((!D !C !B !A)+(!D !C !B A)+(!D !C B !A)+(!D !C B A)+(!D C !B !A)+(!D C !B A)+(!D C B !A)+(!D C B A)), LSE_LINE_FILE_ID=3, LSE_LCOL=13, LSE_RCOL=44, LSE_LLINE=32, LSE_RLINE=32 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(11[2:53])
    defparam I1.init = 16'b0000000011111111;
    
endmodule
//
// Verilog Description of module inverter_U448
//

module inverter_U448 (\notGate[595]_keep , \notGate[596] ) /* synthesis syn_module_defined=1 */ ;
    input \notGate[595]_keep ;
    output \notGate[596] ;
    
    wire \notGate[595]_keep  /* synthesis alspreserve=1 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(25[15:22])
    
    LUT4 I1 (.A(\notGate[595]_keep ), .B(\notGate[595]_keep ), .C(\notGate[595]_keep ), 
         .D(\notGate[595]_keep ), .Z(\notGate[596] )) /* synthesis syn_instantiated=1, lut_function=((!D !C !B !A)+(!D !C !B A)+(!D !C B !A)+(!D !C B A)+(!D C !B !A)+(!D C !B A)+(!D C B !A)+(!D C B A)), LSE_LINE_FILE_ID=3, LSE_LCOL=13, LSE_RCOL=44, LSE_LLINE=32, LSE_RLINE=32 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(11[2:53])
    defparam I1.init = 16'b0000000011111111;
    
endmodule
//
// Verilog Description of module inverter_U449
//

module inverter_U449 (\notGate[594]_keep , \notGate[595] ) /* synthesis syn_module_defined=1 */ ;
    input \notGate[594]_keep ;
    output \notGate[595] ;
    
    wire \notGate[594]_keep  /* synthesis alspreserve=1 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(25[15:22])
    
    LUT4 I1 (.A(\notGate[594]_keep ), .B(\notGate[594]_keep ), .C(\notGate[594]_keep ), 
         .D(\notGate[594]_keep ), .Z(\notGate[595] )) /* synthesis syn_instantiated=1, lut_function=((!D !C !B !A)+(!D !C !B A)+(!D !C B !A)+(!D !C B A)+(!D C !B !A)+(!D C !B A)+(!D C B !A)+(!D C B A)), LSE_LINE_FILE_ID=3, LSE_LCOL=13, LSE_RCOL=44, LSE_LLINE=32, LSE_RLINE=32 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(11[2:53])
    defparam I1.init = 16'b0000000011111111;
    
endmodule
//
// Verilog Description of module inverter_U450
//

module inverter_U450 (\notGate[593]_keep , \notGate[594] ) /* synthesis syn_module_defined=1 */ ;
    input \notGate[593]_keep ;
    output \notGate[594] ;
    
    wire \notGate[593]_keep  /* synthesis alspreserve=1 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(25[15:22])
    
    LUT4 I1 (.A(\notGate[593]_keep ), .B(\notGate[593]_keep ), .C(\notGate[593]_keep ), 
         .D(\notGate[593]_keep ), .Z(\notGate[594] )) /* synthesis syn_instantiated=1, lut_function=((!D !C !B !A)+(!D !C !B A)+(!D !C B !A)+(!D !C B A)+(!D C !B !A)+(!D C !B A)+(!D C B !A)+(!D C B A)), LSE_LINE_FILE_ID=3, LSE_LCOL=13, LSE_RCOL=44, LSE_LLINE=32, LSE_RLINE=32 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(11[2:53])
    defparam I1.init = 16'b0000000011111111;
    
endmodule
//
// Verilog Description of module inverter_U451
//

module inverter_U451 (\notGate[592]_keep , \notGate[593] ) /* synthesis syn_module_defined=1 */ ;
    input \notGate[592]_keep ;
    output \notGate[593] ;
    
    wire \notGate[592]_keep  /* synthesis alspreserve=1 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(25[15:22])
    
    LUT4 I1 (.A(\notGate[592]_keep ), .B(\notGate[592]_keep ), .C(\notGate[592]_keep ), 
         .D(\notGate[592]_keep ), .Z(\notGate[593] )) /* synthesis syn_instantiated=1, lut_function=((!D !C !B !A)+(!D !C !B A)+(!D !C B !A)+(!D !C B A)+(!D C !B !A)+(!D C !B A)+(!D C B !A)+(!D C B A)), LSE_LINE_FILE_ID=3, LSE_LCOL=13, LSE_RCOL=44, LSE_LLINE=32, LSE_RLINE=32 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(11[2:53])
    defparam I1.init = 16'b0000000011111111;
    
endmodule
//
// Verilog Description of module inverter_U452
//

module inverter_U452 (\notGate[591]_keep , \notGate[592] ) /* synthesis syn_module_defined=1 */ ;
    input \notGate[591]_keep ;
    output \notGate[592] ;
    
    wire \notGate[591]_keep  /* synthesis alspreserve=1 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(25[15:22])
    
    LUT4 I1 (.A(\notGate[591]_keep ), .B(\notGate[591]_keep ), .C(\notGate[591]_keep ), 
         .D(\notGate[591]_keep ), .Z(\notGate[592] )) /* synthesis syn_instantiated=1, lut_function=((!D !C !B !A)+(!D !C !B A)+(!D !C B !A)+(!D !C B A)+(!D C !B !A)+(!D C !B A)+(!D C B !A)+(!D C B A)), LSE_LINE_FILE_ID=3, LSE_LCOL=13, LSE_RCOL=44, LSE_LLINE=32, LSE_RLINE=32 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(11[2:53])
    defparam I1.init = 16'b0000000011111111;
    
endmodule
//
// Verilog Description of module inverter_U453
//

module inverter_U453 (\notGate[590]_keep , \notGate[591] ) /* synthesis syn_module_defined=1 */ ;
    input \notGate[590]_keep ;
    output \notGate[591] ;
    
    wire \notGate[590]_keep  /* synthesis alspreserve=1 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(25[15:22])
    
    LUT4 I1 (.A(\notGate[590]_keep ), .B(\notGate[590]_keep ), .C(\notGate[590]_keep ), 
         .D(\notGate[590]_keep ), .Z(\notGate[591] )) /* synthesis syn_instantiated=1, lut_function=((!D !C !B !A)+(!D !C !B A)+(!D !C B !A)+(!D !C B A)+(!D C !B !A)+(!D C !B A)+(!D C B !A)+(!D C B A)), LSE_LINE_FILE_ID=3, LSE_LCOL=13, LSE_RCOL=44, LSE_LLINE=32, LSE_RLINE=32 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(11[2:53])
    defparam I1.init = 16'b0000000011111111;
    
endmodule
//
// Verilog Description of module inverter_U454
//

module inverter_U454 (\notGate[589]_keep , \notGate[590] ) /* synthesis syn_module_defined=1 */ ;
    input \notGate[589]_keep ;
    output \notGate[590] ;
    
    wire \notGate[589]_keep  /* synthesis alspreserve=1 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(25[15:22])
    
    LUT4 I1 (.A(\notGate[589]_keep ), .B(\notGate[589]_keep ), .C(\notGate[589]_keep ), 
         .D(\notGate[589]_keep ), .Z(\notGate[590] )) /* synthesis syn_instantiated=1, lut_function=((!D !C !B !A)+(!D !C !B A)+(!D !C B !A)+(!D !C B A)+(!D C !B !A)+(!D C !B A)+(!D C B !A)+(!D C B A)), LSE_LINE_FILE_ID=3, LSE_LCOL=13, LSE_RCOL=44, LSE_LLINE=32, LSE_RLINE=32 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(11[2:53])
    defparam I1.init = 16'b0000000011111111;
    
endmodule
//
// Verilog Description of module inverter_U455
//

module inverter_U455 (\notGate[57]_keep , \notGate[58] ) /* synthesis syn_module_defined=1 */ ;
    input \notGate[57]_keep ;
    output \notGate[58] ;
    
    wire \notGate[57]_keep  /* synthesis alspreserve=1 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(25[15:22])
    
    LUT4 I1 (.A(\notGate[57]_keep ), .B(\notGate[57]_keep ), .C(\notGate[57]_keep ), 
         .D(\notGate[57]_keep ), .Z(\notGate[58] )) /* synthesis syn_instantiated=1, lut_function=((!D !C !B !A)+(!D !C !B A)+(!D !C B !A)+(!D !C B A)+(!D C !B !A)+(!D C !B A)+(!D C B !A)+(!D C B A)), LSE_LINE_FILE_ID=3, LSE_LCOL=13, LSE_RCOL=44, LSE_LLINE=32, LSE_RLINE=32 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(11[2:53])
    defparam I1.init = 16'b0000000011111111;
    
endmodule
//
// Verilog Description of module inverter_U456
//

module inverter_U456 (\notGate[588]_keep , \notGate[589] ) /* synthesis syn_module_defined=1 */ ;
    input \notGate[588]_keep ;
    output \notGate[589] ;
    
    wire \notGate[588]_keep  /* synthesis alspreserve=1 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(25[15:22])
    
    LUT4 I1 (.A(\notGate[588]_keep ), .B(\notGate[588]_keep ), .C(\notGate[588]_keep ), 
         .D(\notGate[588]_keep ), .Z(\notGate[589] )) /* synthesis syn_instantiated=1, lut_function=((!D !C !B !A)+(!D !C !B A)+(!D !C B !A)+(!D !C B A)+(!D C !B !A)+(!D C !B A)+(!D C B !A)+(!D C B A)), LSE_LINE_FILE_ID=3, LSE_LCOL=13, LSE_RCOL=44, LSE_LLINE=32, LSE_RLINE=32 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(11[2:53])
    defparam I1.init = 16'b0000000011111111;
    
endmodule
//
// Verilog Description of module inverter_U457
//

module inverter_U457 (\notGate[587]_keep , \notGate[588] ) /* synthesis syn_module_defined=1 */ ;
    input \notGate[587]_keep ;
    output \notGate[588] ;
    
    wire \notGate[587]_keep  /* synthesis alspreserve=1 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(25[15:22])
    
    LUT4 I1 (.A(\notGate[587]_keep ), .B(\notGate[587]_keep ), .C(\notGate[587]_keep ), 
         .D(\notGate[587]_keep ), .Z(\notGate[588] )) /* synthesis syn_instantiated=1, lut_function=((!D !C !B !A)+(!D !C !B A)+(!D !C B !A)+(!D !C B A)+(!D C !B !A)+(!D C !B A)+(!D C B !A)+(!D C B A)), LSE_LINE_FILE_ID=3, LSE_LCOL=13, LSE_RCOL=44, LSE_LLINE=32, LSE_RLINE=32 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(11[2:53])
    defparam I1.init = 16'b0000000011111111;
    
endmodule
//
// Verilog Description of module inverter_U458
//

module inverter_U458 (\notGate[586]_keep , \notGate[587] ) /* synthesis syn_module_defined=1 */ ;
    input \notGate[586]_keep ;
    output \notGate[587] ;
    
    wire \notGate[586]_keep  /* synthesis alspreserve=1 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(25[15:22])
    
    LUT4 I1 (.A(\notGate[586]_keep ), .B(\notGate[586]_keep ), .C(\notGate[586]_keep ), 
         .D(\notGate[586]_keep ), .Z(\notGate[587] )) /* synthesis syn_instantiated=1, lut_function=((!D !C !B !A)+(!D !C !B A)+(!D !C B !A)+(!D !C B A)+(!D C !B !A)+(!D C !B A)+(!D C B !A)+(!D C B A)), LSE_LINE_FILE_ID=3, LSE_LCOL=13, LSE_RCOL=44, LSE_LLINE=32, LSE_RLINE=32 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(11[2:53])
    defparam I1.init = 16'b0000000011111111;
    
endmodule
//
// Verilog Description of module inverter_U459
//

module inverter_U459 (\notGate[585]_keep , \notGate[586] ) /* synthesis syn_module_defined=1 */ ;
    input \notGate[585]_keep ;
    output \notGate[586] ;
    
    wire \notGate[585]_keep  /* synthesis alspreserve=1 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(25[15:22])
    
    LUT4 I1 (.A(\notGate[585]_keep ), .B(\notGate[585]_keep ), .C(\notGate[585]_keep ), 
         .D(\notGate[585]_keep ), .Z(\notGate[586] )) /* synthesis syn_instantiated=1, lut_function=((!D !C !B !A)+(!D !C !B A)+(!D !C B !A)+(!D !C B A)+(!D C !B !A)+(!D C !B A)+(!D C B !A)+(!D C B A)), LSE_LINE_FILE_ID=3, LSE_LCOL=13, LSE_RCOL=44, LSE_LLINE=32, LSE_RLINE=32 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(11[2:53])
    defparam I1.init = 16'b0000000011111111;
    
endmodule
//
// Verilog Description of module inverter_U460
//

module inverter_U460 (\notGate[584]_keep , \notGate[585] ) /* synthesis syn_module_defined=1 */ ;
    input \notGate[584]_keep ;
    output \notGate[585] ;
    
    wire \notGate[584]_keep  /* synthesis alspreserve=1 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(25[15:22])
    
    LUT4 I1 (.A(\notGate[584]_keep ), .B(\notGate[584]_keep ), .C(\notGate[584]_keep ), 
         .D(\notGate[584]_keep ), .Z(\notGate[585] )) /* synthesis syn_instantiated=1, lut_function=((!D !C !B !A)+(!D !C !B A)+(!D !C B !A)+(!D !C B A)+(!D C !B !A)+(!D C !B A)+(!D C B !A)+(!D C B A)), LSE_LINE_FILE_ID=3, LSE_LCOL=13, LSE_RCOL=44, LSE_LLINE=32, LSE_RLINE=32 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(11[2:53])
    defparam I1.init = 16'b0000000011111111;
    
endmodule
//
// Verilog Description of module inverter_U461
//

module inverter_U461 (\notGate[583]_keep , \notGate[584] ) /* synthesis syn_module_defined=1 */ ;
    input \notGate[583]_keep ;
    output \notGate[584] ;
    
    wire \notGate[583]_keep  /* synthesis alspreserve=1 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(25[15:22])
    
    LUT4 I1 (.A(\notGate[583]_keep ), .B(\notGate[583]_keep ), .C(\notGate[583]_keep ), 
         .D(\notGate[583]_keep ), .Z(\notGate[584] )) /* synthesis syn_instantiated=1, lut_function=((!D !C !B !A)+(!D !C !B A)+(!D !C B !A)+(!D !C B A)+(!D C !B !A)+(!D C !B A)+(!D C B !A)+(!D C B A)), LSE_LINE_FILE_ID=3, LSE_LCOL=13, LSE_RCOL=44, LSE_LLINE=32, LSE_RLINE=32 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(11[2:53])
    defparam I1.init = 16'b0000000011111111;
    
endmodule
//
// Verilog Description of module inverter_U462
//

module inverter_U462 (\notGate[582]_keep , \notGate[583] ) /* synthesis syn_module_defined=1 */ ;
    input \notGate[582]_keep ;
    output \notGate[583] ;
    
    wire \notGate[582]_keep  /* synthesis alspreserve=1 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(25[15:22])
    
    LUT4 I1 (.A(\notGate[582]_keep ), .B(\notGate[582]_keep ), .C(\notGate[582]_keep ), 
         .D(\notGate[582]_keep ), .Z(\notGate[583] )) /* synthesis syn_instantiated=1, lut_function=((!D !C !B !A)+(!D !C !B A)+(!D !C B !A)+(!D !C B A)+(!D C !B !A)+(!D C !B A)+(!D C B !A)+(!D C B A)), LSE_LINE_FILE_ID=3, LSE_LCOL=13, LSE_RCOL=44, LSE_LLINE=32, LSE_RLINE=32 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(11[2:53])
    defparam I1.init = 16'b0000000011111111;
    
endmodule
//
// Verilog Description of module inverter_U463
//

module inverter_U463 (\notGate[581]_keep , \notGate[582] ) /* synthesis syn_module_defined=1 */ ;
    input \notGate[581]_keep ;
    output \notGate[582] ;
    
    wire \notGate[581]_keep  /* synthesis alspreserve=1 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(25[15:22])
    
    LUT4 I1 (.A(\notGate[581]_keep ), .B(\notGate[581]_keep ), .C(\notGate[581]_keep ), 
         .D(\notGate[581]_keep ), .Z(\notGate[582] )) /* synthesis syn_instantiated=1, lut_function=((!D !C !B !A)+(!D !C !B A)+(!D !C B !A)+(!D !C B A)+(!D C !B !A)+(!D C !B A)+(!D C B !A)+(!D C B A)), LSE_LINE_FILE_ID=3, LSE_LCOL=13, LSE_RCOL=44, LSE_LLINE=32, LSE_RLINE=32 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(11[2:53])
    defparam I1.init = 16'b0000000011111111;
    
endmodule
//
// Verilog Description of module inverter_U464
//

module inverter_U464 (\notGate[580]_keep , \notGate[581] ) /* synthesis syn_module_defined=1 */ ;
    input \notGate[580]_keep ;
    output \notGate[581] ;
    
    wire \notGate[580]_keep  /* synthesis alspreserve=1 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(25[15:22])
    
    LUT4 I1 (.A(\notGate[580]_keep ), .B(\notGate[580]_keep ), .C(\notGate[580]_keep ), 
         .D(\notGate[580]_keep ), .Z(\notGate[581] )) /* synthesis syn_instantiated=1, lut_function=((!D !C !B !A)+(!D !C !B A)+(!D !C B !A)+(!D !C B A)+(!D C !B !A)+(!D C !B A)+(!D C B !A)+(!D C B A)), LSE_LINE_FILE_ID=3, LSE_LCOL=13, LSE_RCOL=44, LSE_LLINE=32, LSE_RLINE=32 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(11[2:53])
    defparam I1.init = 16'b0000000011111111;
    
endmodule
//
// Verilog Description of module inverter_U465
//

module inverter_U465 (\notGate[579]_keep , \notGate[580] ) /* synthesis syn_module_defined=1 */ ;
    input \notGate[579]_keep ;
    output \notGate[580] ;
    
    wire \notGate[579]_keep  /* synthesis alspreserve=1 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(25[15:22])
    
    LUT4 I1 (.A(\notGate[579]_keep ), .B(\notGate[579]_keep ), .C(\notGate[579]_keep ), 
         .D(\notGate[579]_keep ), .Z(\notGate[580] )) /* synthesis syn_instantiated=1, lut_function=((!D !C !B !A)+(!D !C !B A)+(!D !C B !A)+(!D !C B A)+(!D C !B !A)+(!D C !B A)+(!D C B !A)+(!D C B A)), LSE_LINE_FILE_ID=3, LSE_LCOL=13, LSE_RCOL=44, LSE_LLINE=32, LSE_RLINE=32 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(11[2:53])
    defparam I1.init = 16'b0000000011111111;
    
endmodule
//
// Verilog Description of module inverter_U466
//

module inverter_U466 (\notGate[56]_keep , \notGate[57] ) /* synthesis syn_module_defined=1 */ ;
    input \notGate[56]_keep ;
    output \notGate[57] ;
    
    wire \notGate[56]_keep  /* synthesis alspreserve=1 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(25[15:22])
    
    LUT4 I1 (.A(\notGate[56]_keep ), .B(\notGate[56]_keep ), .C(\notGate[56]_keep ), 
         .D(\notGate[56]_keep ), .Z(\notGate[57] )) /* synthesis syn_instantiated=1, lut_function=((!D !C !B !A)+(!D !C !B A)+(!D !C B !A)+(!D !C B A)+(!D C !B !A)+(!D C !B A)+(!D C B !A)+(!D C B A)), LSE_LINE_FILE_ID=3, LSE_LCOL=13, LSE_RCOL=44, LSE_LLINE=32, LSE_RLINE=32 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(11[2:53])
    defparam I1.init = 16'b0000000011111111;
    
endmodule
//
// Verilog Description of module inverter_U467
//

module inverter_U467 (\notGate[578]_keep , \notGate[579] ) /* synthesis syn_module_defined=1 */ ;
    input \notGate[578]_keep ;
    output \notGate[579] ;
    
    wire \notGate[578]_keep  /* synthesis alspreserve=1 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(25[15:22])
    
    LUT4 I1 (.A(\notGate[578]_keep ), .B(\notGate[578]_keep ), .C(\notGate[578]_keep ), 
         .D(\notGate[578]_keep ), .Z(\notGate[579] )) /* synthesis syn_instantiated=1, lut_function=((!D !C !B !A)+(!D !C !B A)+(!D !C B !A)+(!D !C B A)+(!D C !B !A)+(!D C !B A)+(!D C B !A)+(!D C B A)), LSE_LINE_FILE_ID=3, LSE_LCOL=13, LSE_RCOL=44, LSE_LLINE=32, LSE_RLINE=32 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(11[2:53])
    defparam I1.init = 16'b0000000011111111;
    
endmodule
//
// Verilog Description of module inverter_U468
//

module inverter_U468 (\notGate[577]_keep , \notGate[578] ) /* synthesis syn_module_defined=1 */ ;
    input \notGate[577]_keep ;
    output \notGate[578] ;
    
    wire \notGate[577]_keep  /* synthesis alspreserve=1 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(25[15:22])
    
    LUT4 I1 (.A(\notGate[577]_keep ), .B(\notGate[577]_keep ), .C(\notGate[577]_keep ), 
         .D(\notGate[577]_keep ), .Z(\notGate[578] )) /* synthesis syn_instantiated=1, lut_function=((!D !C !B !A)+(!D !C !B A)+(!D !C B !A)+(!D !C B A)+(!D C !B !A)+(!D C !B A)+(!D C B !A)+(!D C B A)), LSE_LINE_FILE_ID=3, LSE_LCOL=13, LSE_RCOL=44, LSE_LLINE=32, LSE_RLINE=32 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(11[2:53])
    defparam I1.init = 16'b0000000011111111;
    
endmodule
//
// Verilog Description of module inverter_U469
//

module inverter_U469 (\notGate[576]_keep , \notGate[577] ) /* synthesis syn_module_defined=1 */ ;
    input \notGate[576]_keep ;
    output \notGate[577] ;
    
    wire \notGate[576]_keep  /* synthesis alspreserve=1 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(25[15:22])
    
    LUT4 I1 (.A(\notGate[576]_keep ), .B(\notGate[576]_keep ), .C(\notGate[576]_keep ), 
         .D(\notGate[576]_keep ), .Z(\notGate[577] )) /* synthesis syn_instantiated=1, lut_function=((!D !C !B !A)+(!D !C !B A)+(!D !C B !A)+(!D !C B A)+(!D C !B !A)+(!D C !B A)+(!D C B !A)+(!D C B A)), LSE_LINE_FILE_ID=3, LSE_LCOL=13, LSE_RCOL=44, LSE_LLINE=32, LSE_RLINE=32 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(11[2:53])
    defparam I1.init = 16'b0000000011111111;
    
endmodule
//
// Verilog Description of module inverter_U470
//

module inverter_U470 (\notGate[575]_keep , \notGate[576] ) /* synthesis syn_module_defined=1 */ ;
    input \notGate[575]_keep ;
    output \notGate[576] ;
    
    wire \notGate[575]_keep  /* synthesis alspreserve=1 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(25[15:22])
    
    LUT4 I1 (.A(\notGate[575]_keep ), .B(\notGate[575]_keep ), .C(\notGate[575]_keep ), 
         .D(\notGate[575]_keep ), .Z(\notGate[576] )) /* synthesis syn_instantiated=1, lut_function=((!D !C !B !A)+(!D !C !B A)+(!D !C B !A)+(!D !C B A)+(!D C !B !A)+(!D C !B A)+(!D C B !A)+(!D C B A)), LSE_LINE_FILE_ID=3, LSE_LCOL=13, LSE_RCOL=44, LSE_LLINE=32, LSE_RLINE=32 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(11[2:53])
    defparam I1.init = 16'b0000000011111111;
    
endmodule
//
// Verilog Description of module inverter_U471
//

module inverter_U471 (\notGate[574]_keep , \notGate[575] ) /* synthesis syn_module_defined=1 */ ;
    input \notGate[574]_keep ;
    output \notGate[575] ;
    
    wire \notGate[574]_keep  /* synthesis alspreserve=1 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(25[15:22])
    
    LUT4 I1 (.A(\notGate[574]_keep ), .B(\notGate[574]_keep ), .C(\notGate[574]_keep ), 
         .D(\notGate[574]_keep ), .Z(\notGate[575] )) /* synthesis syn_instantiated=1, lut_function=((!D !C !B !A)+(!D !C !B A)+(!D !C B !A)+(!D !C B A)+(!D C !B !A)+(!D C !B A)+(!D C B !A)+(!D C B A)), LSE_LINE_FILE_ID=3, LSE_LCOL=13, LSE_RCOL=44, LSE_LLINE=32, LSE_RLINE=32 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(11[2:53])
    defparam I1.init = 16'b0000000011111111;
    
endmodule
//
// Verilog Description of module inverter_U472
//

module inverter_U472 (\notGate[573]_keep , \notGate[574] ) /* synthesis syn_module_defined=1 */ ;
    input \notGate[573]_keep ;
    output \notGate[574] ;
    
    wire \notGate[573]_keep  /* synthesis alspreserve=1 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(25[15:22])
    
    LUT4 I1 (.A(\notGate[573]_keep ), .B(\notGate[573]_keep ), .C(\notGate[573]_keep ), 
         .D(\notGate[573]_keep ), .Z(\notGate[574] )) /* synthesis syn_instantiated=1, lut_function=((!D !C !B !A)+(!D !C !B A)+(!D !C B !A)+(!D !C B A)+(!D C !B !A)+(!D C !B A)+(!D C B !A)+(!D C B A)), LSE_LINE_FILE_ID=3, LSE_LCOL=13, LSE_RCOL=44, LSE_LLINE=32, LSE_RLINE=32 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(11[2:53])
    defparam I1.init = 16'b0000000011111111;
    
endmodule
//
// Verilog Description of module inverter_U473
//

module inverter_U473 (\notGate[572]_keep , \notGate[573] ) /* synthesis syn_module_defined=1 */ ;
    input \notGate[572]_keep ;
    output \notGate[573] ;
    
    wire \notGate[572]_keep  /* synthesis alspreserve=1 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(25[15:22])
    
    LUT4 I1 (.A(\notGate[572]_keep ), .B(\notGate[572]_keep ), .C(\notGate[572]_keep ), 
         .D(\notGate[572]_keep ), .Z(\notGate[573] )) /* synthesis syn_instantiated=1, lut_function=((!D !C !B !A)+(!D !C !B A)+(!D !C B !A)+(!D !C B A)+(!D C !B !A)+(!D C !B A)+(!D C B !A)+(!D C B A)), LSE_LINE_FILE_ID=3, LSE_LCOL=13, LSE_RCOL=44, LSE_LLINE=32, LSE_RLINE=32 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(11[2:53])
    defparam I1.init = 16'b0000000011111111;
    
endmodule
//
// Verilog Description of module inverter_U474
//

module inverter_U474 (\notGate[571]_keep , \notGate[572] ) /* synthesis syn_module_defined=1 */ ;
    input \notGate[571]_keep ;
    output \notGate[572] ;
    
    wire \notGate[571]_keep  /* synthesis alspreserve=1 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(25[15:22])
    
    LUT4 I1 (.A(\notGate[571]_keep ), .B(\notGate[571]_keep ), .C(\notGate[571]_keep ), 
         .D(\notGate[571]_keep ), .Z(\notGate[572] )) /* synthesis syn_instantiated=1, lut_function=((!D !C !B !A)+(!D !C !B A)+(!D !C B !A)+(!D !C B A)+(!D C !B !A)+(!D C !B A)+(!D C B !A)+(!D C B A)), LSE_LINE_FILE_ID=3, LSE_LCOL=13, LSE_RCOL=44, LSE_LLINE=32, LSE_RLINE=32 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(11[2:53])
    defparam I1.init = 16'b0000000011111111;
    
endmodule
//
// Verilog Description of module inverter_U475
//

module inverter_U475 (\notGate[570]_keep , \notGate[571] ) /* synthesis syn_module_defined=1 */ ;
    input \notGate[570]_keep ;
    output \notGate[571] ;
    
    wire \notGate[570]_keep  /* synthesis alspreserve=1 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(25[15:22])
    
    LUT4 I1 (.A(\notGate[570]_keep ), .B(\notGate[570]_keep ), .C(\notGate[570]_keep ), 
         .D(\notGate[570]_keep ), .Z(\notGate[571] )) /* synthesis syn_instantiated=1, lut_function=((!D !C !B !A)+(!D !C !B A)+(!D !C B !A)+(!D !C B A)+(!D C !B !A)+(!D C !B A)+(!D C B !A)+(!D C B A)), LSE_LINE_FILE_ID=3, LSE_LCOL=13, LSE_RCOL=44, LSE_LLINE=32, LSE_RLINE=32 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(11[2:53])
    defparam I1.init = 16'b0000000011111111;
    
endmodule
//
// Verilog Description of module inverter_U476
//

module inverter_U476 (\notGate[569]_keep , \notGate[570] ) /* synthesis syn_module_defined=1 */ ;
    input \notGate[569]_keep ;
    output \notGate[570] ;
    
    wire \notGate[569]_keep  /* synthesis alspreserve=1 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(25[15:22])
    
    LUT4 I1 (.A(\notGate[569]_keep ), .B(\notGate[569]_keep ), .C(\notGate[569]_keep ), 
         .D(\notGate[569]_keep ), .Z(\notGate[570] )) /* synthesis syn_instantiated=1, lut_function=((!D !C !B !A)+(!D !C !B A)+(!D !C B !A)+(!D !C B A)+(!D C !B !A)+(!D C !B A)+(!D C B !A)+(!D C B A)), LSE_LINE_FILE_ID=3, LSE_LCOL=13, LSE_RCOL=44, LSE_LLINE=32, LSE_RLINE=32 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(11[2:53])
    defparam I1.init = 16'b0000000011111111;
    
endmodule
//
// Verilog Description of module inverter_U477
//

module inverter_U477 (\notGate[55]_keep , \notGate[56] ) /* synthesis syn_module_defined=1 */ ;
    input \notGate[55]_keep ;
    output \notGate[56] ;
    
    wire \notGate[55]_keep  /* synthesis alspreserve=1 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(25[15:22])
    
    LUT4 I1 (.A(\notGate[55]_keep ), .B(\notGate[55]_keep ), .C(\notGate[55]_keep ), 
         .D(\notGate[55]_keep ), .Z(\notGate[56] )) /* synthesis syn_instantiated=1, lut_function=((!D !C !B !A)+(!D !C !B A)+(!D !C B !A)+(!D !C B A)+(!D C !B !A)+(!D C !B A)+(!D C B !A)+(!D C B A)), LSE_LINE_FILE_ID=3, LSE_LCOL=13, LSE_RCOL=44, LSE_LLINE=32, LSE_RLINE=32 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(11[2:53])
    defparam I1.init = 16'b0000000011111111;
    
endmodule
//
// Verilog Description of module inverter_U478
//

module inverter_U478 (\notGate[568]_keep , \notGate[569] ) /* synthesis syn_module_defined=1 */ ;
    input \notGate[568]_keep ;
    output \notGate[569] ;
    
    wire \notGate[568]_keep  /* synthesis alspreserve=1 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(25[15:22])
    
    LUT4 I1 (.A(\notGate[568]_keep ), .B(\notGate[568]_keep ), .C(\notGate[568]_keep ), 
         .D(\notGate[568]_keep ), .Z(\notGate[569] )) /* synthesis syn_instantiated=1, lut_function=((!D !C !B !A)+(!D !C !B A)+(!D !C B !A)+(!D !C B A)+(!D C !B !A)+(!D C !B A)+(!D C B !A)+(!D C B A)), LSE_LINE_FILE_ID=3, LSE_LCOL=13, LSE_RCOL=44, LSE_LLINE=32, LSE_RLINE=32 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(11[2:53])
    defparam I1.init = 16'b0000000011111111;
    
endmodule
//
// Verilog Description of module inverter_U479
//

module inverter_U479 (\notGate[567]_keep , \notGate[568] ) /* synthesis syn_module_defined=1 */ ;
    input \notGate[567]_keep ;
    output \notGate[568] ;
    
    wire \notGate[567]_keep  /* synthesis alspreserve=1 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(25[15:22])
    
    LUT4 I1 (.A(\notGate[567]_keep ), .B(\notGate[567]_keep ), .C(\notGate[567]_keep ), 
         .D(\notGate[567]_keep ), .Z(\notGate[568] )) /* synthesis syn_instantiated=1, lut_function=((!D !C !B !A)+(!D !C !B A)+(!D !C B !A)+(!D !C B A)+(!D C !B !A)+(!D C !B A)+(!D C B !A)+(!D C B A)), LSE_LINE_FILE_ID=3, LSE_LCOL=13, LSE_RCOL=44, LSE_LLINE=32, LSE_RLINE=32 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(11[2:53])
    defparam I1.init = 16'b0000000011111111;
    
endmodule
//
// Verilog Description of module inverter_U480
//

module inverter_U480 (\notGate[566]_keep , \notGate[567] ) /* synthesis syn_module_defined=1 */ ;
    input \notGate[566]_keep ;
    output \notGate[567] ;
    
    wire \notGate[566]_keep  /* synthesis alspreserve=1 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(25[15:22])
    
    LUT4 I1 (.A(\notGate[566]_keep ), .B(\notGate[566]_keep ), .C(\notGate[566]_keep ), 
         .D(\notGate[566]_keep ), .Z(\notGate[567] )) /* synthesis syn_instantiated=1, lut_function=((!D !C !B !A)+(!D !C !B A)+(!D !C B !A)+(!D !C B A)+(!D C !B !A)+(!D C !B A)+(!D C B !A)+(!D C B A)), LSE_LINE_FILE_ID=3, LSE_LCOL=13, LSE_RCOL=44, LSE_LLINE=32, LSE_RLINE=32 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(11[2:53])
    defparam I1.init = 16'b0000000011111111;
    
endmodule
//
// Verilog Description of module inverter_U481
//

module inverter_U481 (\notGate[565]_keep , \notGate[566] ) /* synthesis syn_module_defined=1 */ ;
    input \notGate[565]_keep ;
    output \notGate[566] ;
    
    wire \notGate[565]_keep  /* synthesis alspreserve=1 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(25[15:22])
    
    LUT4 I1 (.A(\notGate[565]_keep ), .B(\notGate[565]_keep ), .C(\notGate[565]_keep ), 
         .D(\notGate[565]_keep ), .Z(\notGate[566] )) /* synthesis syn_instantiated=1, lut_function=((!D !C !B !A)+(!D !C !B A)+(!D !C B !A)+(!D !C B A)+(!D C !B !A)+(!D C !B A)+(!D C B !A)+(!D C B A)), LSE_LINE_FILE_ID=3, LSE_LCOL=13, LSE_RCOL=44, LSE_LLINE=32, LSE_RLINE=32 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(11[2:53])
    defparam I1.init = 16'b0000000011111111;
    
endmodule
//
// Verilog Description of module inverter_U482
//

module inverter_U482 (\notGate[564]_keep , \notGate[565] ) /* synthesis syn_module_defined=1 */ ;
    input \notGate[564]_keep ;
    output \notGate[565] ;
    
    wire \notGate[564]_keep  /* synthesis alspreserve=1 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(25[15:22])
    
    LUT4 I1 (.A(\notGate[564]_keep ), .B(\notGate[564]_keep ), .C(\notGate[564]_keep ), 
         .D(\notGate[564]_keep ), .Z(\notGate[565] )) /* synthesis syn_instantiated=1, lut_function=((!D !C !B !A)+(!D !C !B A)+(!D !C B !A)+(!D !C B A)+(!D C !B !A)+(!D C !B A)+(!D C B !A)+(!D C B A)), LSE_LINE_FILE_ID=3, LSE_LCOL=13, LSE_RCOL=44, LSE_LLINE=32, LSE_RLINE=32 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(11[2:53])
    defparam I1.init = 16'b0000000011111111;
    
endmodule
//
// Verilog Description of module inverter_U483
//

module inverter_U483 (\notGate[563]_keep , \notGate[564] ) /* synthesis syn_module_defined=1 */ ;
    input \notGate[563]_keep ;
    output \notGate[564] ;
    
    wire \notGate[563]_keep  /* synthesis alspreserve=1 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(25[15:22])
    
    LUT4 I1 (.A(\notGate[563]_keep ), .B(\notGate[563]_keep ), .C(\notGate[563]_keep ), 
         .D(\notGate[563]_keep ), .Z(\notGate[564] )) /* synthesis syn_instantiated=1, lut_function=((!D !C !B !A)+(!D !C !B A)+(!D !C B !A)+(!D !C B A)+(!D C !B !A)+(!D C !B A)+(!D C B !A)+(!D C B A)), LSE_LINE_FILE_ID=3, LSE_LCOL=13, LSE_RCOL=44, LSE_LLINE=32, LSE_RLINE=32 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(11[2:53])
    defparam I1.init = 16'b0000000011111111;
    
endmodule
//
// Verilog Description of module inverter_U484
//

module inverter_U484 (\notGate[562]_keep , \notGate[563] ) /* synthesis syn_module_defined=1 */ ;
    input \notGate[562]_keep ;
    output \notGate[563] ;
    
    wire \notGate[562]_keep  /* synthesis alspreserve=1 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(25[15:22])
    
    LUT4 I1 (.A(\notGate[562]_keep ), .B(\notGate[562]_keep ), .C(\notGate[562]_keep ), 
         .D(\notGate[562]_keep ), .Z(\notGate[563] )) /* synthesis syn_instantiated=1, lut_function=((!D !C !B !A)+(!D !C !B A)+(!D !C B !A)+(!D !C B A)+(!D C !B !A)+(!D C !B A)+(!D C B !A)+(!D C B A)), LSE_LINE_FILE_ID=3, LSE_LCOL=13, LSE_RCOL=44, LSE_LLINE=32, LSE_RLINE=32 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(11[2:53])
    defparam I1.init = 16'b0000000011111111;
    
endmodule
//
// Verilog Description of module inverter_U485
//

module inverter_U485 (\notGate[561]_keep , \notGate[562] ) /* synthesis syn_module_defined=1 */ ;
    input \notGate[561]_keep ;
    output \notGate[562] ;
    
    wire \notGate[561]_keep  /* synthesis alspreserve=1 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(25[15:22])
    
    LUT4 I1 (.A(\notGate[561]_keep ), .B(\notGate[561]_keep ), .C(\notGate[561]_keep ), 
         .D(\notGate[561]_keep ), .Z(\notGate[562] )) /* synthesis syn_instantiated=1, lut_function=((!D !C !B !A)+(!D !C !B A)+(!D !C B !A)+(!D !C B A)+(!D C !B !A)+(!D C !B A)+(!D C B !A)+(!D C B A)), LSE_LINE_FILE_ID=3, LSE_LCOL=13, LSE_RCOL=44, LSE_LLINE=32, LSE_RLINE=32 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(11[2:53])
    defparam I1.init = 16'b0000000011111111;
    
endmodule
//
// Verilog Description of module inverter_U486
//

module inverter_U486 (\notGate[560]_keep , \notGate[561] ) /* synthesis syn_module_defined=1 */ ;
    input \notGate[560]_keep ;
    output \notGate[561] ;
    
    wire \notGate[560]_keep  /* synthesis alspreserve=1 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(25[15:22])
    
    LUT4 I1 (.A(\notGate[560]_keep ), .B(\notGate[560]_keep ), .C(\notGate[560]_keep ), 
         .D(\notGate[560]_keep ), .Z(\notGate[561] )) /* synthesis syn_instantiated=1, lut_function=((!D !C !B !A)+(!D !C !B A)+(!D !C B !A)+(!D !C B A)+(!D C !B !A)+(!D C !B A)+(!D C B !A)+(!D C B A)), LSE_LINE_FILE_ID=3, LSE_LCOL=13, LSE_RCOL=44, LSE_LLINE=32, LSE_RLINE=32 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(11[2:53])
    defparam I1.init = 16'b0000000011111111;
    
endmodule
//
// Verilog Description of module inverter_U487
//

module inverter_U487 (\notGate[559]_keep , \notGate[560] ) /* synthesis syn_module_defined=1 */ ;
    input \notGate[559]_keep ;
    output \notGate[560] ;
    
    wire \notGate[559]_keep  /* synthesis alspreserve=1 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(25[15:22])
    
    LUT4 I1 (.A(\notGate[559]_keep ), .B(\notGate[559]_keep ), .C(\notGate[559]_keep ), 
         .D(\notGate[559]_keep ), .Z(\notGate[560] )) /* synthesis syn_instantiated=1, lut_function=((!D !C !B !A)+(!D !C !B A)+(!D !C B !A)+(!D !C B A)+(!D C !B !A)+(!D C !B A)+(!D C B !A)+(!D C B A)), LSE_LINE_FILE_ID=3, LSE_LCOL=13, LSE_RCOL=44, LSE_LLINE=32, LSE_RLINE=32 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(11[2:53])
    defparam I1.init = 16'b0000000011111111;
    
endmodule
//
// Verilog Description of module inverter_U488
//

module inverter_U488 (\notGate[54]_keep , \notGate[55] ) /* synthesis syn_module_defined=1 */ ;
    input \notGate[54]_keep ;
    output \notGate[55] ;
    
    wire \notGate[54]_keep  /* synthesis alspreserve=1 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(25[15:22])
    
    LUT4 I1 (.A(\notGate[54]_keep ), .B(\notGate[54]_keep ), .C(\notGate[54]_keep ), 
         .D(\notGate[54]_keep ), .Z(\notGate[55] )) /* synthesis syn_instantiated=1, lut_function=((!D !C !B !A)+(!D !C !B A)+(!D !C B !A)+(!D !C B A)+(!D C !B !A)+(!D C !B A)+(!D C B !A)+(!D C B A)), LSE_LINE_FILE_ID=3, LSE_LCOL=13, LSE_RCOL=44, LSE_LLINE=32, LSE_RLINE=32 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(11[2:53])
    defparam I1.init = 16'b0000000011111111;
    
endmodule
//
// Verilog Description of module inverter_U489
//

module inverter_U489 (\notGate[558]_keep , \notGate[559] ) /* synthesis syn_module_defined=1 */ ;
    input \notGate[558]_keep ;
    output \notGate[559] ;
    
    wire \notGate[558]_keep  /* synthesis alspreserve=1 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(25[15:22])
    
    LUT4 I1 (.A(\notGate[558]_keep ), .B(\notGate[558]_keep ), .C(\notGate[558]_keep ), 
         .D(\notGate[558]_keep ), .Z(\notGate[559] )) /* synthesis syn_instantiated=1, lut_function=((!D !C !B !A)+(!D !C !B A)+(!D !C B !A)+(!D !C B A)+(!D C !B !A)+(!D C !B A)+(!D C B !A)+(!D C B A)), LSE_LINE_FILE_ID=3, LSE_LCOL=13, LSE_RCOL=44, LSE_LLINE=32, LSE_RLINE=32 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(11[2:53])
    defparam I1.init = 16'b0000000011111111;
    
endmodule
//
// Verilog Description of module inverter_U490
//

module inverter_U490 (\notGate[557]_keep , \notGate[558] ) /* synthesis syn_module_defined=1 */ ;
    input \notGate[557]_keep ;
    output \notGate[558] ;
    
    wire \notGate[557]_keep  /* synthesis alspreserve=1 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(25[15:22])
    
    LUT4 I1 (.A(\notGate[557]_keep ), .B(\notGate[557]_keep ), .C(\notGate[557]_keep ), 
         .D(\notGate[557]_keep ), .Z(\notGate[558] )) /* synthesis syn_instantiated=1, lut_function=((!D !C !B !A)+(!D !C !B A)+(!D !C B !A)+(!D !C B A)+(!D C !B !A)+(!D C !B A)+(!D C B !A)+(!D C B A)), LSE_LINE_FILE_ID=3, LSE_LCOL=13, LSE_RCOL=44, LSE_LLINE=32, LSE_RLINE=32 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(11[2:53])
    defparam I1.init = 16'b0000000011111111;
    
endmodule
//
// Verilog Description of module inverter_U491
//

module inverter_U491 (\notGate[556]_keep , \notGate[557] ) /* synthesis syn_module_defined=1 */ ;
    input \notGate[556]_keep ;
    output \notGate[557] ;
    
    wire \notGate[556]_keep  /* synthesis alspreserve=1 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(25[15:22])
    
    LUT4 I1 (.A(\notGate[556]_keep ), .B(\notGate[556]_keep ), .C(\notGate[556]_keep ), 
         .D(\notGate[556]_keep ), .Z(\notGate[557] )) /* synthesis syn_instantiated=1, lut_function=((!D !C !B !A)+(!D !C !B A)+(!D !C B !A)+(!D !C B A)+(!D C !B !A)+(!D C !B A)+(!D C B !A)+(!D C B A)), LSE_LINE_FILE_ID=3, LSE_LCOL=13, LSE_RCOL=44, LSE_LLINE=32, LSE_RLINE=32 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(11[2:53])
    defparam I1.init = 16'b0000000011111111;
    
endmodule
//
// Verilog Description of module inverter_U492
//

module inverter_U492 (\notGate[555]_keep , \notGate[556] ) /* synthesis syn_module_defined=1 */ ;
    input \notGate[555]_keep ;
    output \notGate[556] ;
    
    wire \notGate[555]_keep  /* synthesis alspreserve=1 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(25[15:22])
    
    LUT4 I1 (.A(\notGate[555]_keep ), .B(\notGate[555]_keep ), .C(\notGate[555]_keep ), 
         .D(\notGate[555]_keep ), .Z(\notGate[556] )) /* synthesis syn_instantiated=1, lut_function=((!D !C !B !A)+(!D !C !B A)+(!D !C B !A)+(!D !C B A)+(!D C !B !A)+(!D C !B A)+(!D C B !A)+(!D C B A)), LSE_LINE_FILE_ID=3, LSE_LCOL=13, LSE_RCOL=44, LSE_LLINE=32, LSE_RLINE=32 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(11[2:53])
    defparam I1.init = 16'b0000000011111111;
    
endmodule
//
// Verilog Description of module inverter_U493
//

module inverter_U493 (\notGate[554]_keep , \notGate[555] ) /* synthesis syn_module_defined=1 */ ;
    input \notGate[554]_keep ;
    output \notGate[555] ;
    
    wire \notGate[554]_keep  /* synthesis alspreserve=1 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(25[15:22])
    
    LUT4 I1 (.A(\notGate[554]_keep ), .B(\notGate[554]_keep ), .C(\notGate[554]_keep ), 
         .D(\notGate[554]_keep ), .Z(\notGate[555] )) /* synthesis syn_instantiated=1, lut_function=((!D !C !B !A)+(!D !C !B A)+(!D !C B !A)+(!D !C B A)+(!D C !B !A)+(!D C !B A)+(!D C B !A)+(!D C B A)), LSE_LINE_FILE_ID=3, LSE_LCOL=13, LSE_RCOL=44, LSE_LLINE=32, LSE_RLINE=32 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(11[2:53])
    defparam I1.init = 16'b0000000011111111;
    
endmodule
//
// Verilog Description of module inverter_U494
//

module inverter_U494 (\notGate[553]_keep , \notGate[554] ) /* synthesis syn_module_defined=1 */ ;
    input \notGate[553]_keep ;
    output \notGate[554] ;
    
    wire \notGate[553]_keep  /* synthesis alspreserve=1 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(25[15:22])
    
    LUT4 I1 (.A(\notGate[553]_keep ), .B(\notGate[553]_keep ), .C(\notGate[553]_keep ), 
         .D(\notGate[553]_keep ), .Z(\notGate[554] )) /* synthesis syn_instantiated=1, lut_function=((!D !C !B !A)+(!D !C !B A)+(!D !C B !A)+(!D !C B A)+(!D C !B !A)+(!D C !B A)+(!D C B !A)+(!D C B A)), LSE_LINE_FILE_ID=3, LSE_LCOL=13, LSE_RCOL=44, LSE_LLINE=32, LSE_RLINE=32 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(11[2:53])
    defparam I1.init = 16'b0000000011111111;
    
endmodule
//
// Verilog Description of module inverter_U495
//

module inverter_U495 (\notGate[552]_keep , \notGate[553] ) /* synthesis syn_module_defined=1 */ ;
    input \notGate[552]_keep ;
    output \notGate[553] ;
    
    wire \notGate[552]_keep  /* synthesis alspreserve=1 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(25[15:22])
    
    LUT4 I1 (.A(\notGate[552]_keep ), .B(\notGate[552]_keep ), .C(\notGate[552]_keep ), 
         .D(\notGate[552]_keep ), .Z(\notGate[553] )) /* synthesis syn_instantiated=1, lut_function=((!D !C !B !A)+(!D !C !B A)+(!D !C B !A)+(!D !C B A)+(!D C !B !A)+(!D C !B A)+(!D C B !A)+(!D C B A)), LSE_LINE_FILE_ID=3, LSE_LCOL=13, LSE_RCOL=44, LSE_LLINE=32, LSE_RLINE=32 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(11[2:53])
    defparam I1.init = 16'b0000000011111111;
    
endmodule
//
// Verilog Description of module inverter_U496
//

module inverter_U496 (\notGate[551]_keep , \notGate[552] ) /* synthesis syn_module_defined=1 */ ;
    input \notGate[551]_keep ;
    output \notGate[552] ;
    
    wire \notGate[551]_keep  /* synthesis alspreserve=1 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(25[15:22])
    
    LUT4 I1 (.A(\notGate[551]_keep ), .B(\notGate[551]_keep ), .C(\notGate[551]_keep ), 
         .D(\notGate[551]_keep ), .Z(\notGate[552] )) /* synthesis syn_instantiated=1, lut_function=((!D !C !B !A)+(!D !C !B A)+(!D !C B !A)+(!D !C B A)+(!D C !B !A)+(!D C !B A)+(!D C B !A)+(!D C B A)), LSE_LINE_FILE_ID=3, LSE_LCOL=13, LSE_RCOL=44, LSE_LLINE=32, LSE_RLINE=32 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(11[2:53])
    defparam I1.init = 16'b0000000011111111;
    
endmodule
//
// Verilog Description of module inverter_U497
//

module inverter_U497 (\notGate[550]_keep , \notGate[551] ) /* synthesis syn_module_defined=1 */ ;
    input \notGate[550]_keep ;
    output \notGate[551] ;
    
    wire \notGate[550]_keep  /* synthesis alspreserve=1 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(25[15:22])
    
    LUT4 I1 (.A(\notGate[550]_keep ), .B(\notGate[550]_keep ), .C(\notGate[550]_keep ), 
         .D(\notGate[550]_keep ), .Z(\notGate[551] )) /* synthesis syn_instantiated=1, lut_function=((!D !C !B !A)+(!D !C !B A)+(!D !C B !A)+(!D !C B A)+(!D C !B !A)+(!D C !B A)+(!D C B !A)+(!D C B A)), LSE_LINE_FILE_ID=3, LSE_LCOL=13, LSE_RCOL=44, LSE_LLINE=32, LSE_RLINE=32 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(11[2:53])
    defparam I1.init = 16'b0000000011111111;
    
endmodule
//
// Verilog Description of module inverter_U498
//

module inverter_U498 (\notGate[549]_keep , \notGate[550] ) /* synthesis syn_module_defined=1 */ ;
    input \notGate[549]_keep ;
    output \notGate[550] ;
    
    wire \notGate[549]_keep  /* synthesis alspreserve=1 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(25[15:22])
    
    LUT4 I1 (.A(\notGate[549]_keep ), .B(\notGate[549]_keep ), .C(\notGate[549]_keep ), 
         .D(\notGate[549]_keep ), .Z(\notGate[550] )) /* synthesis syn_instantiated=1, lut_function=((!D !C !B !A)+(!D !C !B A)+(!D !C B !A)+(!D !C B A)+(!D C !B !A)+(!D C !B A)+(!D C B !A)+(!D C B A)), LSE_LINE_FILE_ID=3, LSE_LCOL=13, LSE_RCOL=44, LSE_LLINE=32, LSE_RLINE=32 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(11[2:53])
    defparam I1.init = 16'b0000000011111111;
    
endmodule
//
// Verilog Description of module inverter_U499
//

module inverter_U499 (\notGate[53]_keep , \notGate[54] ) /* synthesis syn_module_defined=1 */ ;
    input \notGate[53]_keep ;
    output \notGate[54] ;
    
    wire \notGate[53]_keep  /* synthesis alspreserve=1 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(25[15:22])
    
    LUT4 I1 (.A(\notGate[53]_keep ), .B(\notGate[53]_keep ), .C(\notGate[53]_keep ), 
         .D(\notGate[53]_keep ), .Z(\notGate[54] )) /* synthesis syn_instantiated=1, lut_function=((!D !C !B !A)+(!D !C !B A)+(!D !C B !A)+(!D !C B A)+(!D C !B !A)+(!D C !B A)+(!D C B !A)+(!D C B A)), LSE_LINE_FILE_ID=3, LSE_LCOL=13, LSE_RCOL=44, LSE_LLINE=32, LSE_RLINE=32 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(11[2:53])
    defparam I1.init = 16'b0000000011111111;
    
endmodule
//
// Verilog Description of module inverter_U500
//

module inverter_U500 (\notGate[548]_keep , \notGate[549] ) /* synthesis syn_module_defined=1 */ ;
    input \notGate[548]_keep ;
    output \notGate[549] ;
    
    wire \notGate[548]_keep  /* synthesis alspreserve=1 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(25[15:22])
    
    LUT4 I1 (.A(\notGate[548]_keep ), .B(\notGate[548]_keep ), .C(\notGate[548]_keep ), 
         .D(\notGate[548]_keep ), .Z(\notGate[549] )) /* synthesis syn_instantiated=1, lut_function=((!D !C !B !A)+(!D !C !B A)+(!D !C B !A)+(!D !C B A)+(!D C !B !A)+(!D C !B A)+(!D C B !A)+(!D C B A)), LSE_LINE_FILE_ID=3, LSE_LCOL=13, LSE_RCOL=44, LSE_LLINE=32, LSE_RLINE=32 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(11[2:53])
    defparam I1.init = 16'b0000000011111111;
    
endmodule
//
// Verilog Description of module inverter_U501
//

module inverter_U501 (\notGate[547]_keep , \notGate[548] ) /* synthesis syn_module_defined=1 */ ;
    input \notGate[547]_keep ;
    output \notGate[548] ;
    
    wire \notGate[547]_keep  /* synthesis alspreserve=1 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(25[15:22])
    
    LUT4 I1 (.A(\notGate[547]_keep ), .B(\notGate[547]_keep ), .C(\notGate[547]_keep ), 
         .D(\notGate[547]_keep ), .Z(\notGate[548] )) /* synthesis syn_instantiated=1, lut_function=((!D !C !B !A)+(!D !C !B A)+(!D !C B !A)+(!D !C B A)+(!D C !B !A)+(!D C !B A)+(!D C B !A)+(!D C B A)), LSE_LINE_FILE_ID=3, LSE_LCOL=13, LSE_RCOL=44, LSE_LLINE=32, LSE_RLINE=32 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(11[2:53])
    defparam I1.init = 16'b0000000011111111;
    
endmodule
//
// Verilog Description of module inverter_U502
//

module inverter_U502 (\notGate[546]_keep , \notGate[547] ) /* synthesis syn_module_defined=1 */ ;
    input \notGate[546]_keep ;
    output \notGate[547] ;
    
    wire \notGate[546]_keep  /* synthesis alspreserve=1 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(25[15:22])
    
    LUT4 I1 (.A(\notGate[546]_keep ), .B(\notGate[546]_keep ), .C(\notGate[546]_keep ), 
         .D(\notGate[546]_keep ), .Z(\notGate[547] )) /* synthesis syn_instantiated=1, lut_function=((!D !C !B !A)+(!D !C !B A)+(!D !C B !A)+(!D !C B A)+(!D C !B !A)+(!D C !B A)+(!D C B !A)+(!D C B A)), LSE_LINE_FILE_ID=3, LSE_LCOL=13, LSE_RCOL=44, LSE_LLINE=32, LSE_RLINE=32 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(11[2:53])
    defparam I1.init = 16'b0000000011111111;
    
endmodule
//
// Verilog Description of module inverter_U503
//

module inverter_U503 (\notGate[545]_keep , \notGate[546] ) /* synthesis syn_module_defined=1 */ ;
    input \notGate[545]_keep ;
    output \notGate[546] ;
    
    wire \notGate[545]_keep  /* synthesis alspreserve=1 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(25[15:22])
    
    LUT4 I1 (.A(\notGate[545]_keep ), .B(\notGate[545]_keep ), .C(\notGate[545]_keep ), 
         .D(\notGate[545]_keep ), .Z(\notGate[546] )) /* synthesis syn_instantiated=1, lut_function=((!D !C !B !A)+(!D !C !B A)+(!D !C B !A)+(!D !C B A)+(!D C !B !A)+(!D C !B A)+(!D C B !A)+(!D C B A)), LSE_LINE_FILE_ID=3, LSE_LCOL=13, LSE_RCOL=44, LSE_LLINE=32, LSE_RLINE=32 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(11[2:53])
    defparam I1.init = 16'b0000000011111111;
    
endmodule
//
// Verilog Description of module inverter_U504
//

module inverter_U504 (\notGate[544]_keep , \notGate[545] ) /* synthesis syn_module_defined=1 */ ;
    input \notGate[544]_keep ;
    output \notGate[545] ;
    
    wire \notGate[544]_keep  /* synthesis alspreserve=1 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(25[15:22])
    
    LUT4 I1 (.A(\notGate[544]_keep ), .B(\notGate[544]_keep ), .C(\notGate[544]_keep ), 
         .D(\notGate[544]_keep ), .Z(\notGate[545] )) /* synthesis syn_instantiated=1, lut_function=((!D !C !B !A)+(!D !C !B A)+(!D !C B !A)+(!D !C B A)+(!D C !B !A)+(!D C !B A)+(!D C B !A)+(!D C B A)), LSE_LINE_FILE_ID=3, LSE_LCOL=13, LSE_RCOL=44, LSE_LLINE=32, LSE_RLINE=32 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(11[2:53])
    defparam I1.init = 16'b0000000011111111;
    
endmodule
//
// Verilog Description of module inverter_U505
//

module inverter_U505 (\notGate[543]_keep , \notGate[544] ) /* synthesis syn_module_defined=1 */ ;
    input \notGate[543]_keep ;
    output \notGate[544] ;
    
    wire \notGate[543]_keep  /* synthesis alspreserve=1 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(25[15:22])
    
    LUT4 I1 (.A(\notGate[543]_keep ), .B(\notGate[543]_keep ), .C(\notGate[543]_keep ), 
         .D(\notGate[543]_keep ), .Z(\notGate[544] )) /* synthesis syn_instantiated=1, lut_function=((!D !C !B !A)+(!D !C !B A)+(!D !C B !A)+(!D !C B A)+(!D C !B !A)+(!D C !B A)+(!D C B !A)+(!D C B A)), LSE_LINE_FILE_ID=3, LSE_LCOL=13, LSE_RCOL=44, LSE_LLINE=32, LSE_RLINE=32 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(11[2:53])
    defparam I1.init = 16'b0000000011111111;
    
endmodule
//
// Verilog Description of module inverter_U506
//

module inverter_U506 (\notGate[542]_keep , \notGate[543] ) /* synthesis syn_module_defined=1 */ ;
    input \notGate[542]_keep ;
    output \notGate[543] ;
    
    wire \notGate[542]_keep  /* synthesis alspreserve=1 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(25[15:22])
    
    LUT4 I1 (.A(\notGate[542]_keep ), .B(\notGate[542]_keep ), .C(\notGate[542]_keep ), 
         .D(\notGate[542]_keep ), .Z(\notGate[543] )) /* synthesis syn_instantiated=1, lut_function=((!D !C !B !A)+(!D !C !B A)+(!D !C B !A)+(!D !C B A)+(!D C !B !A)+(!D C !B A)+(!D C B !A)+(!D C B A)), LSE_LINE_FILE_ID=3, LSE_LCOL=13, LSE_RCOL=44, LSE_LLINE=32, LSE_RLINE=32 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(11[2:53])
    defparam I1.init = 16'b0000000011111111;
    
endmodule
//
// Verilog Description of module inverter_U507
//

module inverter_U507 (\notGate[541]_keep , \notGate[542] ) /* synthesis syn_module_defined=1 */ ;
    input \notGate[541]_keep ;
    output \notGate[542] ;
    
    wire \notGate[541]_keep  /* synthesis alspreserve=1 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(25[15:22])
    
    LUT4 I1 (.A(\notGate[541]_keep ), .B(\notGate[541]_keep ), .C(\notGate[541]_keep ), 
         .D(\notGate[541]_keep ), .Z(\notGate[542] )) /* synthesis syn_instantiated=1, lut_function=((!D !C !B !A)+(!D !C !B A)+(!D !C B !A)+(!D !C B A)+(!D C !B !A)+(!D C !B A)+(!D C B !A)+(!D C B A)), LSE_LINE_FILE_ID=3, LSE_LCOL=13, LSE_RCOL=44, LSE_LLINE=32, LSE_RLINE=32 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(11[2:53])
    defparam I1.init = 16'b0000000011111111;
    
endmodule
//
// Verilog Description of module inverter_U508
//

module inverter_U508 (\notGate[540]_keep , \notGate[541] ) /* synthesis syn_module_defined=1 */ ;
    input \notGate[540]_keep ;
    output \notGate[541] ;
    
    wire \notGate[540]_keep  /* synthesis alspreserve=1 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(25[15:22])
    
    LUT4 I1 (.A(\notGate[540]_keep ), .B(\notGate[540]_keep ), .C(\notGate[540]_keep ), 
         .D(\notGate[540]_keep ), .Z(\notGate[541] )) /* synthesis syn_instantiated=1, lut_function=((!D !C !B !A)+(!D !C !B A)+(!D !C B !A)+(!D !C B A)+(!D C !B !A)+(!D C !B A)+(!D C B !A)+(!D C B A)), LSE_LINE_FILE_ID=3, LSE_LCOL=13, LSE_RCOL=44, LSE_LLINE=32, LSE_RLINE=32 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(11[2:53])
    defparam I1.init = 16'b0000000011111111;
    
endmodule
//
// Verilog Description of module inverter_U509
//

module inverter_U509 (\notGate[539]_keep , \notGate[540] ) /* synthesis syn_module_defined=1 */ ;
    input \notGate[539]_keep ;
    output \notGate[540] ;
    
    wire \notGate[539]_keep  /* synthesis alspreserve=1 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(25[15:22])
    
    LUT4 I1 (.A(\notGate[539]_keep ), .B(\notGate[539]_keep ), .C(\notGate[539]_keep ), 
         .D(\notGate[539]_keep ), .Z(\notGate[540] )) /* synthesis syn_instantiated=1, lut_function=((!D !C !B !A)+(!D !C !B A)+(!D !C B !A)+(!D !C B A)+(!D C !B !A)+(!D C !B A)+(!D C B !A)+(!D C B A)), LSE_LINE_FILE_ID=3, LSE_LCOL=13, LSE_RCOL=44, LSE_LLINE=32, LSE_RLINE=32 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(11[2:53])
    defparam I1.init = 16'b0000000011111111;
    
endmodule
//
// Verilog Description of module inverter_U510
//

module inverter_U510 (\notGate[52]_keep , \notGate[53] ) /* synthesis syn_module_defined=1 */ ;
    input \notGate[52]_keep ;
    output \notGate[53] ;
    
    wire \notGate[52]_keep  /* synthesis alspreserve=1 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(25[15:22])
    
    LUT4 I1 (.A(\notGate[52]_keep ), .B(\notGate[52]_keep ), .C(\notGate[52]_keep ), 
         .D(\notGate[52]_keep ), .Z(\notGate[53] )) /* synthesis syn_instantiated=1, lut_function=((!D !C !B !A)+(!D !C !B A)+(!D !C B !A)+(!D !C B A)+(!D C !B !A)+(!D C !B A)+(!D C B !A)+(!D C B A)), LSE_LINE_FILE_ID=3, LSE_LCOL=13, LSE_RCOL=44, LSE_LLINE=32, LSE_RLINE=32 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(11[2:53])
    defparam I1.init = 16'b0000000011111111;
    
endmodule
//
// Verilog Description of module inverter_U511
//

module inverter_U511 (\notGate[538]_keep , \notGate[539] ) /* synthesis syn_module_defined=1 */ ;
    input \notGate[538]_keep ;
    output \notGate[539] ;
    
    wire \notGate[538]_keep  /* synthesis alspreserve=1 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(25[15:22])
    
    LUT4 I1 (.A(\notGate[538]_keep ), .B(\notGate[538]_keep ), .C(\notGate[538]_keep ), 
         .D(\notGate[538]_keep ), .Z(\notGate[539] )) /* synthesis syn_instantiated=1, lut_function=((!D !C !B !A)+(!D !C !B A)+(!D !C B !A)+(!D !C B A)+(!D C !B !A)+(!D C !B A)+(!D C B !A)+(!D C B A)), LSE_LINE_FILE_ID=3, LSE_LCOL=13, LSE_RCOL=44, LSE_LLINE=32, LSE_RLINE=32 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(11[2:53])
    defparam I1.init = 16'b0000000011111111;
    
endmodule
//
// Verilog Description of module inverter_U512
//

module inverter_U512 (\notGate[537]_keep , \notGate[538] ) /* synthesis syn_module_defined=1 */ ;
    input \notGate[537]_keep ;
    output \notGate[538] ;
    
    wire \notGate[537]_keep  /* synthesis alspreserve=1 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(25[15:22])
    
    LUT4 I1 (.A(\notGate[537]_keep ), .B(\notGate[537]_keep ), .C(\notGate[537]_keep ), 
         .D(\notGate[537]_keep ), .Z(\notGate[538] )) /* synthesis syn_instantiated=1, lut_function=((!D !C !B !A)+(!D !C !B A)+(!D !C B !A)+(!D !C B A)+(!D C !B !A)+(!D C !B A)+(!D C B !A)+(!D C B A)), LSE_LINE_FILE_ID=3, LSE_LCOL=13, LSE_RCOL=44, LSE_LLINE=32, LSE_RLINE=32 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(11[2:53])
    defparam I1.init = 16'b0000000011111111;
    
endmodule
//
// Verilog Description of module inverter_U513
//

module inverter_U513 (\notGate[536]_keep , \notGate[537] ) /* synthesis syn_module_defined=1 */ ;
    input \notGate[536]_keep ;
    output \notGate[537] ;
    
    wire \notGate[536]_keep  /* synthesis alspreserve=1 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(25[15:22])
    
    LUT4 I1 (.A(\notGate[536]_keep ), .B(\notGate[536]_keep ), .C(\notGate[536]_keep ), 
         .D(\notGate[536]_keep ), .Z(\notGate[537] )) /* synthesis syn_instantiated=1, lut_function=((!D !C !B !A)+(!D !C !B A)+(!D !C B !A)+(!D !C B A)+(!D C !B !A)+(!D C !B A)+(!D C B !A)+(!D C B A)), LSE_LINE_FILE_ID=3, LSE_LCOL=13, LSE_RCOL=44, LSE_LLINE=32, LSE_RLINE=32 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(11[2:53])
    defparam I1.init = 16'b0000000011111111;
    
endmodule
//
// Verilog Description of module inverter_U514
//

module inverter_U514 (\notGate[535]_keep , \notGate[536] ) /* synthesis syn_module_defined=1 */ ;
    input \notGate[535]_keep ;
    output \notGate[536] ;
    
    wire \notGate[535]_keep  /* synthesis alspreserve=1 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(25[15:22])
    
    LUT4 I1 (.A(\notGate[535]_keep ), .B(\notGate[535]_keep ), .C(\notGate[535]_keep ), 
         .D(\notGate[535]_keep ), .Z(\notGate[536] )) /* synthesis syn_instantiated=1, lut_function=((!D !C !B !A)+(!D !C !B A)+(!D !C B !A)+(!D !C B A)+(!D C !B !A)+(!D C !B A)+(!D C B !A)+(!D C B A)), LSE_LINE_FILE_ID=3, LSE_LCOL=13, LSE_RCOL=44, LSE_LLINE=32, LSE_RLINE=32 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(11[2:53])
    defparam I1.init = 16'b0000000011111111;
    
endmodule
//
// Verilog Description of module inverter_U515
//

module inverter_U515 (\notGate[534]_keep , \notGate[535] ) /* synthesis syn_module_defined=1 */ ;
    input \notGate[534]_keep ;
    output \notGate[535] ;
    
    wire \notGate[534]_keep  /* synthesis alspreserve=1 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(25[15:22])
    
    LUT4 I1 (.A(\notGate[534]_keep ), .B(\notGate[534]_keep ), .C(\notGate[534]_keep ), 
         .D(\notGate[534]_keep ), .Z(\notGate[535] )) /* synthesis syn_instantiated=1, lut_function=((!D !C !B !A)+(!D !C !B A)+(!D !C B !A)+(!D !C B A)+(!D C !B !A)+(!D C !B A)+(!D C B !A)+(!D C B A)), LSE_LINE_FILE_ID=3, LSE_LCOL=13, LSE_RCOL=44, LSE_LLINE=32, LSE_RLINE=32 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(11[2:53])
    defparam I1.init = 16'b0000000011111111;
    
endmodule
//
// Verilog Description of module inverter_U516
//

module inverter_U516 (\notGate[533]_keep , \notGate[534] ) /* synthesis syn_module_defined=1 */ ;
    input \notGate[533]_keep ;
    output \notGate[534] ;
    
    wire \notGate[533]_keep  /* synthesis alspreserve=1 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(25[15:22])
    
    LUT4 I1 (.A(\notGate[533]_keep ), .B(\notGate[533]_keep ), .C(\notGate[533]_keep ), 
         .D(\notGate[533]_keep ), .Z(\notGate[534] )) /* synthesis syn_instantiated=1, lut_function=((!D !C !B !A)+(!D !C !B A)+(!D !C B !A)+(!D !C B A)+(!D C !B !A)+(!D C !B A)+(!D C B !A)+(!D C B A)), LSE_LINE_FILE_ID=3, LSE_LCOL=13, LSE_RCOL=44, LSE_LLINE=32, LSE_RLINE=32 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(11[2:53])
    defparam I1.init = 16'b0000000011111111;
    
endmodule
//
// Verilog Description of module inverter_U517
//

module inverter_U517 (\notGate[532]_keep , \notGate[533] ) /* synthesis syn_module_defined=1 */ ;
    input \notGate[532]_keep ;
    output \notGate[533] ;
    
    wire \notGate[532]_keep  /* synthesis alspreserve=1 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(25[15:22])
    
    LUT4 I1 (.A(\notGate[532]_keep ), .B(\notGate[532]_keep ), .C(\notGate[532]_keep ), 
         .D(\notGate[532]_keep ), .Z(\notGate[533] )) /* synthesis syn_instantiated=1, lut_function=((!D !C !B !A)+(!D !C !B A)+(!D !C B !A)+(!D !C B A)+(!D C !B !A)+(!D C !B A)+(!D C B !A)+(!D C B A)), LSE_LINE_FILE_ID=3, LSE_LCOL=13, LSE_RCOL=44, LSE_LLINE=32, LSE_RLINE=32 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(11[2:53])
    defparam I1.init = 16'b0000000011111111;
    
endmodule
//
// Verilog Description of module inverter_U518
//

module inverter_U518 (\notGate[531]_keep , \notGate[532] ) /* synthesis syn_module_defined=1 */ ;
    input \notGate[531]_keep ;
    output \notGate[532] ;
    
    wire \notGate[531]_keep  /* synthesis alspreserve=1 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(25[15:22])
    
    LUT4 I1 (.A(\notGate[531]_keep ), .B(\notGate[531]_keep ), .C(\notGate[531]_keep ), 
         .D(\notGate[531]_keep ), .Z(\notGate[532] )) /* synthesis syn_instantiated=1, lut_function=((!D !C !B !A)+(!D !C !B A)+(!D !C B !A)+(!D !C B A)+(!D C !B !A)+(!D C !B A)+(!D C B !A)+(!D C B A)), LSE_LINE_FILE_ID=3, LSE_LCOL=13, LSE_RCOL=44, LSE_LLINE=32, LSE_RLINE=32 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(11[2:53])
    defparam I1.init = 16'b0000000011111111;
    
endmodule
//
// Verilog Description of module inverter_U519
//

module inverter_U519 (\notGate[530]_keep , \notGate[531] ) /* synthesis syn_module_defined=1 */ ;
    input \notGate[530]_keep ;
    output \notGate[531] ;
    
    wire \notGate[530]_keep  /* synthesis alspreserve=1 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(25[15:22])
    
    LUT4 I1 (.A(\notGate[530]_keep ), .B(\notGate[530]_keep ), .C(\notGate[530]_keep ), 
         .D(\notGate[530]_keep ), .Z(\notGate[531] )) /* synthesis syn_instantiated=1, lut_function=((!D !C !B !A)+(!D !C !B A)+(!D !C B !A)+(!D !C B A)+(!D C !B !A)+(!D C !B A)+(!D C B !A)+(!D C B A)), LSE_LINE_FILE_ID=3, LSE_LCOL=13, LSE_RCOL=44, LSE_LLINE=32, LSE_RLINE=32 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(11[2:53])
    defparam I1.init = 16'b0000000011111111;
    
endmodule
//
// Verilog Description of module inverter_U520
//

module inverter_U520 (\notGate[529]_keep , \notGate[530] ) /* synthesis syn_module_defined=1 */ ;
    input \notGate[529]_keep ;
    output \notGate[530] ;
    
    wire \notGate[529]_keep  /* synthesis alspreserve=1 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(25[15:22])
    
    LUT4 I1 (.A(\notGate[529]_keep ), .B(\notGate[529]_keep ), .C(\notGate[529]_keep ), 
         .D(\notGate[529]_keep ), .Z(\notGate[530] )) /* synthesis syn_instantiated=1, lut_function=((!D !C !B !A)+(!D !C !B A)+(!D !C B !A)+(!D !C B A)+(!D C !B !A)+(!D C !B A)+(!D C B !A)+(!D C B A)), LSE_LINE_FILE_ID=3, LSE_LCOL=13, LSE_RCOL=44, LSE_LLINE=32, LSE_RLINE=32 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(11[2:53])
    defparam I1.init = 16'b0000000011111111;
    
endmodule
//
// Verilog Description of module inverter_U521
//

module inverter_U521 (\notGate[51]_keep , \notGate[52] ) /* synthesis syn_module_defined=1 */ ;
    input \notGate[51]_keep ;
    output \notGate[52] ;
    
    wire \notGate[51]_keep  /* synthesis alspreserve=1 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(25[15:22])
    
    LUT4 I1 (.A(\notGate[51]_keep ), .B(\notGate[51]_keep ), .C(\notGate[51]_keep ), 
         .D(\notGate[51]_keep ), .Z(\notGate[52] )) /* synthesis syn_instantiated=1, lut_function=((!D !C !B !A)+(!D !C !B A)+(!D !C B !A)+(!D !C B A)+(!D C !B !A)+(!D C !B A)+(!D C B !A)+(!D C B A)), LSE_LINE_FILE_ID=3, LSE_LCOL=13, LSE_RCOL=44, LSE_LLINE=32, LSE_RLINE=32 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(11[2:53])
    defparam I1.init = 16'b0000000011111111;
    
endmodule
//
// Verilog Description of module inverter_U522
//

module inverter_U522 (\notGate[528]_keep , \notGate[529] ) /* synthesis syn_module_defined=1 */ ;
    input \notGate[528]_keep ;
    output \notGate[529] ;
    
    wire \notGate[528]_keep  /* synthesis alspreserve=1 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(25[15:22])
    
    LUT4 I1 (.A(\notGate[528]_keep ), .B(\notGate[528]_keep ), .C(\notGate[528]_keep ), 
         .D(\notGate[528]_keep ), .Z(\notGate[529] )) /* synthesis syn_instantiated=1, lut_function=((!D !C !B !A)+(!D !C !B A)+(!D !C B !A)+(!D !C B A)+(!D C !B !A)+(!D C !B A)+(!D C B !A)+(!D C B A)), LSE_LINE_FILE_ID=3, LSE_LCOL=13, LSE_RCOL=44, LSE_LLINE=32, LSE_RLINE=32 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(11[2:53])
    defparam I1.init = 16'b0000000011111111;
    
endmodule
//
// Verilog Description of module inverter_U523
//

module inverter_U523 (\notGate[527]_keep , \notGate[528] ) /* synthesis syn_module_defined=1 */ ;
    input \notGate[527]_keep ;
    output \notGate[528] ;
    
    wire \notGate[527]_keep  /* synthesis alspreserve=1 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(25[15:22])
    
    LUT4 I1 (.A(\notGate[527]_keep ), .B(\notGate[527]_keep ), .C(\notGate[527]_keep ), 
         .D(\notGate[527]_keep ), .Z(\notGate[528] )) /* synthesis syn_instantiated=1, lut_function=((!D !C !B !A)+(!D !C !B A)+(!D !C B !A)+(!D !C B A)+(!D C !B !A)+(!D C !B A)+(!D C B !A)+(!D C B A)), LSE_LINE_FILE_ID=3, LSE_LCOL=13, LSE_RCOL=44, LSE_LLINE=32, LSE_RLINE=32 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(11[2:53])
    defparam I1.init = 16'b0000000011111111;
    
endmodule
//
// Verilog Description of module inverter_U524
//

module inverter_U524 (\notGate[526]_keep , \notGate[527] ) /* synthesis syn_module_defined=1 */ ;
    input \notGate[526]_keep ;
    output \notGate[527] ;
    
    wire \notGate[526]_keep  /* synthesis alspreserve=1 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(25[15:22])
    
    LUT4 I1 (.A(\notGate[526]_keep ), .B(\notGate[526]_keep ), .C(\notGate[526]_keep ), 
         .D(\notGate[526]_keep ), .Z(\notGate[527] )) /* synthesis syn_instantiated=1, lut_function=((!D !C !B !A)+(!D !C !B A)+(!D !C B !A)+(!D !C B A)+(!D C !B !A)+(!D C !B A)+(!D C B !A)+(!D C B A)), LSE_LINE_FILE_ID=3, LSE_LCOL=13, LSE_RCOL=44, LSE_LLINE=32, LSE_RLINE=32 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(11[2:53])
    defparam I1.init = 16'b0000000011111111;
    
endmodule
//
// Verilog Description of module inverter_U525
//

module inverter_U525 (\notGate[525]_keep , \notGate[526] ) /* synthesis syn_module_defined=1 */ ;
    input \notGate[525]_keep ;
    output \notGate[526] ;
    
    wire \notGate[525]_keep  /* synthesis alspreserve=1 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(25[15:22])
    
    LUT4 I1 (.A(\notGate[525]_keep ), .B(\notGate[525]_keep ), .C(\notGate[525]_keep ), 
         .D(\notGate[525]_keep ), .Z(\notGate[526] )) /* synthesis syn_instantiated=1, lut_function=((!D !C !B !A)+(!D !C !B A)+(!D !C B !A)+(!D !C B A)+(!D C !B !A)+(!D C !B A)+(!D C B !A)+(!D C B A)), LSE_LINE_FILE_ID=3, LSE_LCOL=13, LSE_RCOL=44, LSE_LLINE=32, LSE_RLINE=32 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(11[2:53])
    defparam I1.init = 16'b0000000011111111;
    
endmodule
//
// Verilog Description of module inverter_U526
//

module inverter_U526 (\notGate[524]_keep , \notGate[525] ) /* synthesis syn_module_defined=1 */ ;
    input \notGate[524]_keep ;
    output \notGate[525] ;
    
    wire \notGate[524]_keep  /* synthesis alspreserve=1 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(25[15:22])
    
    LUT4 I1 (.A(\notGate[524]_keep ), .B(\notGate[524]_keep ), .C(\notGate[524]_keep ), 
         .D(\notGate[524]_keep ), .Z(\notGate[525] )) /* synthesis syn_instantiated=1, lut_function=((!D !C !B !A)+(!D !C !B A)+(!D !C B !A)+(!D !C B A)+(!D C !B !A)+(!D C !B A)+(!D C B !A)+(!D C B A)), LSE_LINE_FILE_ID=3, LSE_LCOL=13, LSE_RCOL=44, LSE_LLINE=32, LSE_RLINE=32 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(11[2:53])
    defparam I1.init = 16'b0000000011111111;
    
endmodule
//
// Verilog Description of module inverter_U527
//

module inverter_U527 (\notGate[523]_keep , \notGate[524] ) /* synthesis syn_module_defined=1 */ ;
    input \notGate[523]_keep ;
    output \notGate[524] ;
    
    wire \notGate[523]_keep  /* synthesis alspreserve=1 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(25[15:22])
    
    LUT4 I1 (.A(\notGate[523]_keep ), .B(\notGate[523]_keep ), .C(\notGate[523]_keep ), 
         .D(\notGate[523]_keep ), .Z(\notGate[524] )) /* synthesis syn_instantiated=1, lut_function=((!D !C !B !A)+(!D !C !B A)+(!D !C B !A)+(!D !C B A)+(!D C !B !A)+(!D C !B A)+(!D C B !A)+(!D C B A)), LSE_LINE_FILE_ID=3, LSE_LCOL=13, LSE_RCOL=44, LSE_LLINE=32, LSE_RLINE=32 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(11[2:53])
    defparam I1.init = 16'b0000000011111111;
    
endmodule
//
// Verilog Description of module inverter_U528
//

module inverter_U528 (\notGate[522]_keep , \notGate[523] ) /* synthesis syn_module_defined=1 */ ;
    input \notGate[522]_keep ;
    output \notGate[523] ;
    
    wire \notGate[522]_keep  /* synthesis alspreserve=1 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(25[15:22])
    
    LUT4 I1 (.A(\notGate[522]_keep ), .B(\notGate[522]_keep ), .C(\notGate[522]_keep ), 
         .D(\notGate[522]_keep ), .Z(\notGate[523] )) /* synthesis syn_instantiated=1, lut_function=((!D !C !B !A)+(!D !C !B A)+(!D !C B !A)+(!D !C B A)+(!D C !B !A)+(!D C !B A)+(!D C B !A)+(!D C B A)), LSE_LINE_FILE_ID=3, LSE_LCOL=13, LSE_RCOL=44, LSE_LLINE=32, LSE_RLINE=32 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(11[2:53])
    defparam I1.init = 16'b0000000011111111;
    
endmodule
//
// Verilog Description of module inverter_U529
//

module inverter_U529 (\notGate[521]_keep , \notGate[522] ) /* synthesis syn_module_defined=1 */ ;
    input \notGate[521]_keep ;
    output \notGate[522] ;
    
    wire \notGate[521]_keep  /* synthesis alspreserve=1 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(25[15:22])
    
    LUT4 I1 (.A(\notGate[521]_keep ), .B(\notGate[521]_keep ), .C(\notGate[521]_keep ), 
         .D(\notGate[521]_keep ), .Z(\notGate[522] )) /* synthesis syn_instantiated=1, lut_function=((!D !C !B !A)+(!D !C !B A)+(!D !C B !A)+(!D !C B A)+(!D C !B !A)+(!D C !B A)+(!D C B !A)+(!D C B A)), LSE_LINE_FILE_ID=3, LSE_LCOL=13, LSE_RCOL=44, LSE_LLINE=32, LSE_RLINE=32 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(11[2:53])
    defparam I1.init = 16'b0000000011111111;
    
endmodule
//
// Verilog Description of module inverter_U530
//

module inverter_U530 (\notGate[520]_keep , \notGate[521] ) /* synthesis syn_module_defined=1 */ ;
    input \notGate[520]_keep ;
    output \notGate[521] ;
    
    wire \notGate[520]_keep  /* synthesis alspreserve=1 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(25[15:22])
    
    LUT4 I1 (.A(\notGate[520]_keep ), .B(\notGate[520]_keep ), .C(\notGate[520]_keep ), 
         .D(\notGate[520]_keep ), .Z(\notGate[521] )) /* synthesis syn_instantiated=1, lut_function=((!D !C !B !A)+(!D !C !B A)+(!D !C B !A)+(!D !C B A)+(!D C !B !A)+(!D C !B A)+(!D C B !A)+(!D C B A)), LSE_LINE_FILE_ID=3, LSE_LCOL=13, LSE_RCOL=44, LSE_LLINE=32, LSE_RLINE=32 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(11[2:53])
    defparam I1.init = 16'b0000000011111111;
    
endmodule
//
// Verilog Description of module inverter_U531
//

module inverter_U531 (\notGate[519]_keep , \notGate[520] ) /* synthesis syn_module_defined=1 */ ;
    input \notGate[519]_keep ;
    output \notGate[520] ;
    
    wire \notGate[519]_keep  /* synthesis alspreserve=1 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(25[15:22])
    
    LUT4 I1 (.A(\notGate[519]_keep ), .B(\notGate[519]_keep ), .C(\notGate[519]_keep ), 
         .D(\notGate[519]_keep ), .Z(\notGate[520] )) /* synthesis syn_instantiated=1, lut_function=((!D !C !B !A)+(!D !C !B A)+(!D !C B !A)+(!D !C B A)+(!D C !B !A)+(!D C !B A)+(!D C B !A)+(!D C B A)), LSE_LINE_FILE_ID=3, LSE_LCOL=13, LSE_RCOL=44, LSE_LLINE=32, LSE_RLINE=32 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(11[2:53])
    defparam I1.init = 16'b0000000011111111;
    
endmodule
//
// Verilog Description of module inverter_U532
//

module inverter_U532 (\notGate[50]_keep , \notGate[51] ) /* synthesis syn_module_defined=1 */ ;
    input \notGate[50]_keep ;
    output \notGate[51] ;
    
    wire \notGate[50]_keep  /* synthesis alspreserve=1 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(25[15:22])
    
    LUT4 I1 (.A(\notGate[50]_keep ), .B(\notGate[50]_keep ), .C(\notGate[50]_keep ), 
         .D(\notGate[50]_keep ), .Z(\notGate[51] )) /* synthesis syn_instantiated=1, lut_function=((!D !C !B !A)+(!D !C !B A)+(!D !C B !A)+(!D !C B A)+(!D C !B !A)+(!D C !B A)+(!D C B !A)+(!D C B A)), LSE_LINE_FILE_ID=3, LSE_LCOL=13, LSE_RCOL=44, LSE_LLINE=32, LSE_RLINE=32 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(11[2:53])
    defparam I1.init = 16'b0000000011111111;
    
endmodule
//
// Verilog Description of module inverter_U533
//

module inverter_U533 (\notGate[518]_keep , \notGate[519] ) /* synthesis syn_module_defined=1 */ ;
    input \notGate[518]_keep ;
    output \notGate[519] ;
    
    wire \notGate[518]_keep  /* synthesis alspreserve=1 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(25[15:22])
    
    LUT4 I1 (.A(\notGate[518]_keep ), .B(\notGate[518]_keep ), .C(\notGate[518]_keep ), 
         .D(\notGate[518]_keep ), .Z(\notGate[519] )) /* synthesis syn_instantiated=1, lut_function=((!D !C !B !A)+(!D !C !B A)+(!D !C B !A)+(!D !C B A)+(!D C !B !A)+(!D C !B A)+(!D C B !A)+(!D C B A)), LSE_LINE_FILE_ID=3, LSE_LCOL=13, LSE_RCOL=44, LSE_LLINE=32, LSE_RLINE=32 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(11[2:53])
    defparam I1.init = 16'b0000000011111111;
    
endmodule
//
// Verilog Description of module inverter_U534
//

module inverter_U534 (\notGate[517]_keep , \notGate[518] ) /* synthesis syn_module_defined=1 */ ;
    input \notGate[517]_keep ;
    output \notGate[518] ;
    
    wire \notGate[517]_keep  /* synthesis alspreserve=1 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(25[15:22])
    
    LUT4 I1 (.A(\notGate[517]_keep ), .B(\notGate[517]_keep ), .C(\notGate[517]_keep ), 
         .D(\notGate[517]_keep ), .Z(\notGate[518] )) /* synthesis syn_instantiated=1, lut_function=((!D !C !B !A)+(!D !C !B A)+(!D !C B !A)+(!D !C B A)+(!D C !B !A)+(!D C !B A)+(!D C B !A)+(!D C B A)), LSE_LINE_FILE_ID=3, LSE_LCOL=13, LSE_RCOL=44, LSE_LLINE=32, LSE_RLINE=32 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(11[2:53])
    defparam I1.init = 16'b0000000011111111;
    
endmodule
//
// Verilog Description of module inverter_U535
//

module inverter_U535 (\notGate[516]_keep , \notGate[517] ) /* synthesis syn_module_defined=1 */ ;
    input \notGate[516]_keep ;
    output \notGate[517] ;
    
    wire \notGate[516]_keep  /* synthesis alspreserve=1 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(25[15:22])
    
    LUT4 I1 (.A(\notGate[516]_keep ), .B(\notGate[516]_keep ), .C(\notGate[516]_keep ), 
         .D(\notGate[516]_keep ), .Z(\notGate[517] )) /* synthesis syn_instantiated=1, lut_function=((!D !C !B !A)+(!D !C !B A)+(!D !C B !A)+(!D !C B A)+(!D C !B !A)+(!D C !B A)+(!D C B !A)+(!D C B A)), LSE_LINE_FILE_ID=3, LSE_LCOL=13, LSE_RCOL=44, LSE_LLINE=32, LSE_RLINE=32 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(11[2:53])
    defparam I1.init = 16'b0000000011111111;
    
endmodule
//
// Verilog Description of module inverter_U536
//

module inverter_U536 (\notGate[515]_keep , \notGate[516] ) /* synthesis syn_module_defined=1 */ ;
    input \notGate[515]_keep ;
    output \notGate[516] ;
    
    wire \notGate[515]_keep  /* synthesis alspreserve=1 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(25[15:22])
    
    LUT4 I1 (.A(\notGate[515]_keep ), .B(\notGate[515]_keep ), .C(\notGate[515]_keep ), 
         .D(\notGate[515]_keep ), .Z(\notGate[516] )) /* synthesis syn_instantiated=1, lut_function=((!D !C !B !A)+(!D !C !B A)+(!D !C B !A)+(!D !C B A)+(!D C !B !A)+(!D C !B A)+(!D C B !A)+(!D C B A)), LSE_LINE_FILE_ID=3, LSE_LCOL=13, LSE_RCOL=44, LSE_LLINE=32, LSE_RLINE=32 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(11[2:53])
    defparam I1.init = 16'b0000000011111111;
    
endmodule
//
// Verilog Description of module inverter_U537
//

module inverter_U537 (\notGate[514]_keep , \notGate[515] ) /* synthesis syn_module_defined=1 */ ;
    input \notGate[514]_keep ;
    output \notGate[515] ;
    
    wire \notGate[514]_keep  /* synthesis alspreserve=1 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(25[15:22])
    
    LUT4 I1 (.A(\notGate[514]_keep ), .B(\notGate[514]_keep ), .C(\notGate[514]_keep ), 
         .D(\notGate[514]_keep ), .Z(\notGate[515] )) /* synthesis syn_instantiated=1, lut_function=((!D !C !B !A)+(!D !C !B A)+(!D !C B !A)+(!D !C B A)+(!D C !B !A)+(!D C !B A)+(!D C B !A)+(!D C B A)), LSE_LINE_FILE_ID=3, LSE_LCOL=13, LSE_RCOL=44, LSE_LLINE=32, LSE_RLINE=32 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(11[2:53])
    defparam I1.init = 16'b0000000011111111;
    
endmodule
//
// Verilog Description of module inverter_U538
//

module inverter_U538 (\notGate[513]_keep , \notGate[514] ) /* synthesis syn_module_defined=1 */ ;
    input \notGate[513]_keep ;
    output \notGate[514] ;
    
    wire \notGate[513]_keep  /* synthesis alspreserve=1 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(25[15:22])
    
    LUT4 I1 (.A(\notGate[513]_keep ), .B(\notGate[513]_keep ), .C(\notGate[513]_keep ), 
         .D(\notGate[513]_keep ), .Z(\notGate[514] )) /* synthesis syn_instantiated=1, lut_function=((!D !C !B !A)+(!D !C !B A)+(!D !C B !A)+(!D !C B A)+(!D C !B !A)+(!D C !B A)+(!D C B !A)+(!D C B A)), LSE_LINE_FILE_ID=3, LSE_LCOL=13, LSE_RCOL=44, LSE_LLINE=32, LSE_RLINE=32 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(11[2:53])
    defparam I1.init = 16'b0000000011111111;
    
endmodule
//
// Verilog Description of module inverter_U539
//

module inverter_U539 (\notGate[512]_keep , \notGate[513] ) /* synthesis syn_module_defined=1 */ ;
    input \notGate[512]_keep ;
    output \notGate[513] ;
    
    wire \notGate[512]_keep  /* synthesis alspreserve=1 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(25[15:22])
    
    LUT4 I1 (.A(\notGate[512]_keep ), .B(\notGate[512]_keep ), .C(\notGate[512]_keep ), 
         .D(\notGate[512]_keep ), .Z(\notGate[513] )) /* synthesis syn_instantiated=1, lut_function=((!D !C !B !A)+(!D !C !B A)+(!D !C B !A)+(!D !C B A)+(!D C !B !A)+(!D C !B A)+(!D C B !A)+(!D C B A)), LSE_LINE_FILE_ID=3, LSE_LCOL=13, LSE_RCOL=44, LSE_LLINE=32, LSE_RLINE=32 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(11[2:53])
    defparam I1.init = 16'b0000000011111111;
    
endmodule
//
// Verilog Description of module inverter_U540
//

module inverter_U540 (\notGate[511]_keep , \notGate[512] ) /* synthesis syn_module_defined=1 */ ;
    input \notGate[511]_keep ;
    output \notGate[512] ;
    
    wire \notGate[511]_keep  /* synthesis alspreserve=1 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(25[15:22])
    
    LUT4 I1 (.A(\notGate[511]_keep ), .B(\notGate[511]_keep ), .C(\notGate[511]_keep ), 
         .D(\notGate[511]_keep ), .Z(\notGate[512] )) /* synthesis syn_instantiated=1, lut_function=((!D !C !B !A)+(!D !C !B A)+(!D !C B !A)+(!D !C B A)+(!D C !B !A)+(!D C !B A)+(!D C B !A)+(!D C B A)), LSE_LINE_FILE_ID=3, LSE_LCOL=13, LSE_RCOL=44, LSE_LLINE=32, LSE_RLINE=32 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(11[2:53])
    defparam I1.init = 16'b0000000011111111;
    
endmodule
//
// Verilog Description of module inverter_U541
//

module inverter_U541 (\notGate[510]_keep , \notGate[511] ) /* synthesis syn_module_defined=1 */ ;
    input \notGate[510]_keep ;
    output \notGate[511] ;
    
    wire \notGate[510]_keep  /* synthesis alspreserve=1 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(25[15:22])
    
    LUT4 I1 (.A(\notGate[510]_keep ), .B(\notGate[510]_keep ), .C(\notGate[510]_keep ), 
         .D(\notGate[510]_keep ), .Z(\notGate[511] )) /* synthesis syn_instantiated=1, lut_function=((!D !C !B !A)+(!D !C !B A)+(!D !C B !A)+(!D !C B A)+(!D C !B !A)+(!D C !B A)+(!D C B !A)+(!D C B A)), LSE_LINE_FILE_ID=3, LSE_LCOL=13, LSE_RCOL=44, LSE_LLINE=32, LSE_RLINE=32 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(11[2:53])
    defparam I1.init = 16'b0000000011111111;
    
endmodule
//
// Verilog Description of module inverter_U542
//

module inverter_U542 (\notGate[509]_keep , \notGate[510] ) /* synthesis syn_module_defined=1 */ ;
    input \notGate[509]_keep ;
    output \notGate[510] ;
    
    wire \notGate[509]_keep  /* synthesis alspreserve=1 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(25[15:22])
    
    LUT4 I1 (.A(\notGate[509]_keep ), .B(\notGate[509]_keep ), .C(\notGate[509]_keep ), 
         .D(\notGate[509]_keep ), .Z(\notGate[510] )) /* synthesis syn_instantiated=1, lut_function=((!D !C !B !A)+(!D !C !B A)+(!D !C B !A)+(!D !C B A)+(!D C !B !A)+(!D C !B A)+(!D C B !A)+(!D C B A)), LSE_LINE_FILE_ID=3, LSE_LCOL=13, LSE_RCOL=44, LSE_LLINE=32, LSE_RLINE=32 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(11[2:53])
    defparam I1.init = 16'b0000000011111111;
    
endmodule
//
// Verilog Description of module inverter_U543
//

module inverter_U543 (\notGate[49]_keep , \notGate[50] ) /* synthesis syn_module_defined=1 */ ;
    input \notGate[49]_keep ;
    output \notGate[50] ;
    
    wire \notGate[49]_keep  /* synthesis alspreserve=1 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(25[15:22])
    
    LUT4 I1 (.A(\notGate[49]_keep ), .B(\notGate[49]_keep ), .C(\notGate[49]_keep ), 
         .D(\notGate[49]_keep ), .Z(\notGate[50] )) /* synthesis syn_instantiated=1, lut_function=((!D !C !B !A)+(!D !C !B A)+(!D !C B !A)+(!D !C B A)+(!D C !B !A)+(!D C !B A)+(!D C B !A)+(!D C B A)), LSE_LINE_FILE_ID=3, LSE_LCOL=13, LSE_RCOL=44, LSE_LLINE=32, LSE_RLINE=32 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(11[2:53])
    defparam I1.init = 16'b0000000011111111;
    
endmodule
//
// Verilog Description of module inverter_U544
//

module inverter_U544 (\notGate[508]_keep , \notGate[509] ) /* synthesis syn_module_defined=1 */ ;
    input \notGate[508]_keep ;
    output \notGate[509] ;
    
    wire \notGate[508]_keep  /* synthesis alspreserve=1 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(25[15:22])
    
    LUT4 I1 (.A(\notGate[508]_keep ), .B(\notGate[508]_keep ), .C(\notGate[508]_keep ), 
         .D(\notGate[508]_keep ), .Z(\notGate[509] )) /* synthesis syn_instantiated=1, lut_function=((!D !C !B !A)+(!D !C !B A)+(!D !C B !A)+(!D !C B A)+(!D C !B !A)+(!D C !B A)+(!D C B !A)+(!D C B A)), LSE_LINE_FILE_ID=3, LSE_LCOL=13, LSE_RCOL=44, LSE_LLINE=32, LSE_RLINE=32 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(11[2:53])
    defparam I1.init = 16'b0000000011111111;
    
endmodule
//
// Verilog Description of module inverter_U545
//

module inverter_U545 (\notGate[507]_keep , \notGate[508] ) /* synthesis syn_module_defined=1 */ ;
    input \notGate[507]_keep ;
    output \notGate[508] ;
    
    wire \notGate[507]_keep  /* synthesis alspreserve=1 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(25[15:22])
    
    LUT4 I1 (.A(\notGate[507]_keep ), .B(\notGate[507]_keep ), .C(\notGate[507]_keep ), 
         .D(\notGate[507]_keep ), .Z(\notGate[508] )) /* synthesis syn_instantiated=1, lut_function=((!D !C !B !A)+(!D !C !B A)+(!D !C B !A)+(!D !C B A)+(!D C !B !A)+(!D C !B A)+(!D C B !A)+(!D C B A)), LSE_LINE_FILE_ID=3, LSE_LCOL=13, LSE_RCOL=44, LSE_LLINE=32, LSE_RLINE=32 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(11[2:53])
    defparam I1.init = 16'b0000000011111111;
    
endmodule
//
// Verilog Description of module inverter_U546
//

module inverter_U546 (\notGate[506]_keep , \notGate[507] ) /* synthesis syn_module_defined=1 */ ;
    input \notGate[506]_keep ;
    output \notGate[507] ;
    
    wire \notGate[506]_keep  /* synthesis alspreserve=1 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(25[15:22])
    
    LUT4 I1 (.A(\notGate[506]_keep ), .B(\notGate[506]_keep ), .C(\notGate[506]_keep ), 
         .D(\notGate[506]_keep ), .Z(\notGate[507] )) /* synthesis syn_instantiated=1, lut_function=((!D !C !B !A)+(!D !C !B A)+(!D !C B !A)+(!D !C B A)+(!D C !B !A)+(!D C !B A)+(!D C B !A)+(!D C B A)), LSE_LINE_FILE_ID=3, LSE_LCOL=13, LSE_RCOL=44, LSE_LLINE=32, LSE_RLINE=32 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(11[2:53])
    defparam I1.init = 16'b0000000011111111;
    
endmodule
//
// Verilog Description of module inverter_U547
//

module inverter_U547 (\notGate[505]_keep , \notGate[506] ) /* synthesis syn_module_defined=1 */ ;
    input \notGate[505]_keep ;
    output \notGate[506] ;
    
    wire \notGate[505]_keep  /* synthesis alspreserve=1 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(25[15:22])
    
    LUT4 I1 (.A(\notGate[505]_keep ), .B(\notGate[505]_keep ), .C(\notGate[505]_keep ), 
         .D(\notGate[505]_keep ), .Z(\notGate[506] )) /* synthesis syn_instantiated=1, lut_function=((!D !C !B !A)+(!D !C !B A)+(!D !C B !A)+(!D !C B A)+(!D C !B !A)+(!D C !B A)+(!D C B !A)+(!D C B A)), LSE_LINE_FILE_ID=3, LSE_LCOL=13, LSE_RCOL=44, LSE_LLINE=32, LSE_RLINE=32 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(11[2:53])
    defparam I1.init = 16'b0000000011111111;
    
endmodule
//
// Verilog Description of module inverter_U548
//

module inverter_U548 (\notGate[504]_keep , \notGate[505] ) /* synthesis syn_module_defined=1 */ ;
    input \notGate[504]_keep ;
    output \notGate[505] ;
    
    wire \notGate[504]_keep  /* synthesis alspreserve=1 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(25[15:22])
    
    LUT4 I1 (.A(\notGate[504]_keep ), .B(\notGate[504]_keep ), .C(\notGate[504]_keep ), 
         .D(\notGate[504]_keep ), .Z(\notGate[505] )) /* synthesis syn_instantiated=1, lut_function=((!D !C !B !A)+(!D !C !B A)+(!D !C B !A)+(!D !C B A)+(!D C !B !A)+(!D C !B A)+(!D C B !A)+(!D C B A)), LSE_LINE_FILE_ID=3, LSE_LCOL=13, LSE_RCOL=44, LSE_LLINE=32, LSE_RLINE=32 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(11[2:53])
    defparam I1.init = 16'b0000000011111111;
    
endmodule
//
// Verilog Description of module inverter_U549
//

module inverter_U549 (\notGate[503]_keep , \notGate[504] ) /* synthesis syn_module_defined=1 */ ;
    input \notGate[503]_keep ;
    output \notGate[504] ;
    
    wire \notGate[503]_keep  /* synthesis alspreserve=1 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(25[15:22])
    
    LUT4 I1 (.A(\notGate[503]_keep ), .B(\notGate[503]_keep ), .C(\notGate[503]_keep ), 
         .D(\notGate[503]_keep ), .Z(\notGate[504] )) /* synthesis syn_instantiated=1, lut_function=((!D !C !B !A)+(!D !C !B A)+(!D !C B !A)+(!D !C B A)+(!D C !B !A)+(!D C !B A)+(!D C B !A)+(!D C B A)), LSE_LINE_FILE_ID=3, LSE_LCOL=13, LSE_RCOL=44, LSE_LLINE=32, LSE_RLINE=32 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(11[2:53])
    defparam I1.init = 16'b0000000011111111;
    
endmodule
//
// Verilog Description of module inverter_U550
//

module inverter_U550 (\notGate[502]_keep , \notGate[503] ) /* synthesis syn_module_defined=1 */ ;
    input \notGate[502]_keep ;
    output \notGate[503] ;
    
    wire \notGate[502]_keep  /* synthesis alspreserve=1 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(25[15:22])
    
    LUT4 I1 (.A(\notGate[502]_keep ), .B(\notGate[502]_keep ), .C(\notGate[502]_keep ), 
         .D(\notGate[502]_keep ), .Z(\notGate[503] )) /* synthesis syn_instantiated=1, lut_function=((!D !C !B !A)+(!D !C !B A)+(!D !C B !A)+(!D !C B A)+(!D C !B !A)+(!D C !B A)+(!D C B !A)+(!D C B A)), LSE_LINE_FILE_ID=3, LSE_LCOL=13, LSE_RCOL=44, LSE_LLINE=32, LSE_RLINE=32 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(11[2:53])
    defparam I1.init = 16'b0000000011111111;
    
endmodule
//
// Verilog Description of module inverter_U551
//

module inverter_U551 (\notGate[501]_keep , \notGate[502] ) /* synthesis syn_module_defined=1 */ ;
    input \notGate[501]_keep ;
    output \notGate[502] ;
    
    wire \notGate[501]_keep  /* synthesis alspreserve=1 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(25[15:22])
    
    LUT4 I1 (.A(\notGate[501]_keep ), .B(\notGate[501]_keep ), .C(\notGate[501]_keep ), 
         .D(\notGate[501]_keep ), .Z(\notGate[502] )) /* synthesis syn_instantiated=1, lut_function=((!D !C !B !A)+(!D !C !B A)+(!D !C B !A)+(!D !C B A)+(!D C !B !A)+(!D C !B A)+(!D C B !A)+(!D C B A)), LSE_LINE_FILE_ID=3, LSE_LCOL=13, LSE_RCOL=44, LSE_LLINE=32, LSE_RLINE=32 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(11[2:53])
    defparam I1.init = 16'b0000000011111111;
    
endmodule
//
// Verilog Description of module inverter_U552
//

module inverter_U552 (\notGate[500]_keep , \notGate[501] ) /* synthesis syn_module_defined=1 */ ;
    input \notGate[500]_keep ;
    output \notGate[501] ;
    
    wire \notGate[500]_keep  /* synthesis alspreserve=1 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(25[15:22])
    
    LUT4 I1 (.A(\notGate[500]_keep ), .B(\notGate[500]_keep ), .C(\notGate[500]_keep ), 
         .D(\notGate[500]_keep ), .Z(\notGate[501] )) /* synthesis syn_instantiated=1, lut_function=((!D !C !B !A)+(!D !C !B A)+(!D !C B !A)+(!D !C B A)+(!D C !B !A)+(!D C !B A)+(!D C B !A)+(!D C B A)), LSE_LINE_FILE_ID=3, LSE_LCOL=13, LSE_RCOL=44, LSE_LLINE=32, LSE_RLINE=32 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(11[2:53])
    defparam I1.init = 16'b0000000011111111;
    
endmodule
//
// Verilog Description of module inverter_U553
//

module inverter_U553 (\notGate[499]_keep , \notGate[500] ) /* synthesis syn_module_defined=1 */ ;
    input \notGate[499]_keep ;
    output \notGate[500] ;
    
    wire \notGate[499]_keep  /* synthesis alspreserve=1 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(25[15:22])
    
    LUT4 I1 (.A(\notGate[499]_keep ), .B(\notGate[499]_keep ), .C(\notGate[499]_keep ), 
         .D(\notGate[499]_keep ), .Z(\notGate[500] )) /* synthesis syn_instantiated=1, lut_function=((!D !C !B !A)+(!D !C !B A)+(!D !C B !A)+(!D !C B A)+(!D C !B !A)+(!D C !B A)+(!D C B !A)+(!D C B A)), LSE_LINE_FILE_ID=3, LSE_LCOL=13, LSE_RCOL=44, LSE_LLINE=32, LSE_RLINE=32 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(11[2:53])
    defparam I1.init = 16'b0000000011111111;
    
endmodule
//
// Verilog Description of module inverter_U554
//

module inverter_U554 (\notGate[3]_keep , \notGate[4] ) /* synthesis syn_module_defined=1 */ ;
    input \notGate[3]_keep ;
    output \notGate[4] ;
    
    wire \notGate[3]_keep  /* synthesis alspreserve=1 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(25[15:22])
    
    LUT4 I1 (.A(\notGate[3]_keep ), .B(\notGate[3]_keep ), .C(\notGate[3]_keep ), 
         .D(\notGate[3]_keep ), .Z(\notGate[4] )) /* synthesis syn_instantiated=1, lut_function=((!D !C !B !A)+(!D !C !B A)+(!D !C B !A)+(!D !C B A)+(!D C !B !A)+(!D C !B A)+(!D C B !A)+(!D C B A)), LSE_LINE_FILE_ID=3, LSE_LCOL=13, LSE_RCOL=44, LSE_LLINE=32, LSE_RLINE=32 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(11[2:53])
    defparam I1.init = 16'b0000000011111111;
    
endmodule
//
// Verilog Description of module inverter_U555
//

module inverter_U555 (\notGate[48]_keep , \notGate[49] ) /* synthesis syn_module_defined=1 */ ;
    input \notGate[48]_keep ;
    output \notGate[49] ;
    
    wire \notGate[48]_keep  /* synthesis alspreserve=1 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(25[15:22])
    
    LUT4 I1 (.A(\notGate[48]_keep ), .B(\notGate[48]_keep ), .C(\notGate[48]_keep ), 
         .D(\notGate[48]_keep ), .Z(\notGate[49] )) /* synthesis syn_instantiated=1, lut_function=((!D !C !B !A)+(!D !C !B A)+(!D !C B !A)+(!D !C B A)+(!D C !B !A)+(!D C !B A)+(!D C B !A)+(!D C B A)), LSE_LINE_FILE_ID=3, LSE_LCOL=13, LSE_RCOL=44, LSE_LLINE=32, LSE_RLINE=32 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(11[2:53])
    defparam I1.init = 16'b0000000011111111;
    
endmodule
//
// Verilog Description of module inverter_U556
//

module inverter_U556 (\notGate[498]_keep , \notGate[499] ) /* synthesis syn_module_defined=1 */ ;
    input \notGate[498]_keep ;
    output \notGate[499] ;
    
    wire \notGate[498]_keep  /* synthesis alspreserve=1 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(25[15:22])
    
    LUT4 I1 (.A(\notGate[498]_keep ), .B(\notGate[498]_keep ), .C(\notGate[498]_keep ), 
         .D(\notGate[498]_keep ), .Z(\notGate[499] )) /* synthesis syn_instantiated=1, lut_function=((!D !C !B !A)+(!D !C !B A)+(!D !C B !A)+(!D !C B A)+(!D C !B !A)+(!D C !B A)+(!D C B !A)+(!D C B A)), LSE_LINE_FILE_ID=3, LSE_LCOL=13, LSE_RCOL=44, LSE_LLINE=32, LSE_RLINE=32 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(11[2:53])
    defparam I1.init = 16'b0000000011111111;
    
endmodule
//
// Verilog Description of module inverter_U557
//

module inverter_U557 (\notGate[497]_keep , \notGate[498] ) /* synthesis syn_module_defined=1 */ ;
    input \notGate[497]_keep ;
    output \notGate[498] ;
    
    wire \notGate[497]_keep  /* synthesis alspreserve=1 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(25[15:22])
    
    LUT4 I1 (.A(\notGate[497]_keep ), .B(\notGate[497]_keep ), .C(\notGate[497]_keep ), 
         .D(\notGate[497]_keep ), .Z(\notGate[498] )) /* synthesis syn_instantiated=1, lut_function=((!D !C !B !A)+(!D !C !B A)+(!D !C B !A)+(!D !C B A)+(!D C !B !A)+(!D C !B A)+(!D C B !A)+(!D C B A)), LSE_LINE_FILE_ID=3, LSE_LCOL=13, LSE_RCOL=44, LSE_LLINE=32, LSE_RLINE=32 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(11[2:53])
    defparam I1.init = 16'b0000000011111111;
    
endmodule
//
// Verilog Description of module inverter_U558
//

module inverter_U558 (\notGate[496]_keep , \notGate[497] ) /* synthesis syn_module_defined=1 */ ;
    input \notGate[496]_keep ;
    output \notGate[497] ;
    
    wire \notGate[496]_keep  /* synthesis alspreserve=1 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(25[15:22])
    
    LUT4 I1 (.A(\notGate[496]_keep ), .B(\notGate[496]_keep ), .C(\notGate[496]_keep ), 
         .D(\notGate[496]_keep ), .Z(\notGate[497] )) /* synthesis syn_instantiated=1, lut_function=((!D !C !B !A)+(!D !C !B A)+(!D !C B !A)+(!D !C B A)+(!D C !B !A)+(!D C !B A)+(!D C B !A)+(!D C B A)), LSE_LINE_FILE_ID=3, LSE_LCOL=13, LSE_RCOL=44, LSE_LLINE=32, LSE_RLINE=32 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(11[2:53])
    defparam I1.init = 16'b0000000011111111;
    
endmodule
//
// Verilog Description of module inverter_U559
//

module inverter_U559 (\notGate[495]_keep , \notGate[496] ) /* synthesis syn_module_defined=1 */ ;
    input \notGate[495]_keep ;
    output \notGate[496] ;
    
    wire \notGate[495]_keep  /* synthesis alspreserve=1 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(25[15:22])
    
    LUT4 I1 (.A(\notGate[495]_keep ), .B(\notGate[495]_keep ), .C(\notGate[495]_keep ), 
         .D(\notGate[495]_keep ), .Z(\notGate[496] )) /* synthesis syn_instantiated=1, lut_function=((!D !C !B !A)+(!D !C !B A)+(!D !C B !A)+(!D !C B A)+(!D C !B !A)+(!D C !B A)+(!D C B !A)+(!D C B A)), LSE_LINE_FILE_ID=3, LSE_LCOL=13, LSE_RCOL=44, LSE_LLINE=32, LSE_RLINE=32 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(11[2:53])
    defparam I1.init = 16'b0000000011111111;
    
endmodule
//
// Verilog Description of module inverter_U560
//

module inverter_U560 (\notGate[494]_keep , \notGate[495] ) /* synthesis syn_module_defined=1 */ ;
    input \notGate[494]_keep ;
    output \notGate[495] ;
    
    wire \notGate[494]_keep  /* synthesis alspreserve=1 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(25[15:22])
    
    LUT4 I1 (.A(\notGate[494]_keep ), .B(\notGate[494]_keep ), .C(\notGate[494]_keep ), 
         .D(\notGate[494]_keep ), .Z(\notGate[495] )) /* synthesis syn_instantiated=1, lut_function=((!D !C !B !A)+(!D !C !B A)+(!D !C B !A)+(!D !C B A)+(!D C !B !A)+(!D C !B A)+(!D C B !A)+(!D C B A)), LSE_LINE_FILE_ID=3, LSE_LCOL=13, LSE_RCOL=44, LSE_LLINE=32, LSE_RLINE=32 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(11[2:53])
    defparam I1.init = 16'b0000000011111111;
    
endmodule
//
// Verilog Description of module inverter_U561
//

module inverter_U561 (\notGate[493]_keep , \notGate[494] ) /* synthesis syn_module_defined=1 */ ;
    input \notGate[493]_keep ;
    output \notGate[494] ;
    
    wire \notGate[493]_keep  /* synthesis alspreserve=1 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(25[15:22])
    
    LUT4 I1 (.A(\notGate[493]_keep ), .B(\notGate[493]_keep ), .C(\notGate[493]_keep ), 
         .D(\notGate[493]_keep ), .Z(\notGate[494] )) /* synthesis syn_instantiated=1, lut_function=((!D !C !B !A)+(!D !C !B A)+(!D !C B !A)+(!D !C B A)+(!D C !B !A)+(!D C !B A)+(!D C B !A)+(!D C B A)), LSE_LINE_FILE_ID=3, LSE_LCOL=13, LSE_RCOL=44, LSE_LLINE=32, LSE_RLINE=32 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(11[2:53])
    defparam I1.init = 16'b0000000011111111;
    
endmodule
//
// Verilog Description of module inverter_U562
//

module inverter_U562 (\notGate[492]_keep , \notGate[493] ) /* synthesis syn_module_defined=1 */ ;
    input \notGate[492]_keep ;
    output \notGate[493] ;
    
    wire \notGate[492]_keep  /* synthesis alspreserve=1 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(25[15:22])
    
    LUT4 I1 (.A(\notGate[492]_keep ), .B(\notGate[492]_keep ), .C(\notGate[492]_keep ), 
         .D(\notGate[492]_keep ), .Z(\notGate[493] )) /* synthesis syn_instantiated=1, lut_function=((!D !C !B !A)+(!D !C !B A)+(!D !C B !A)+(!D !C B A)+(!D C !B !A)+(!D C !B A)+(!D C B !A)+(!D C B A)), LSE_LINE_FILE_ID=3, LSE_LCOL=13, LSE_RCOL=44, LSE_LLINE=32, LSE_RLINE=32 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(11[2:53])
    defparam I1.init = 16'b0000000011111111;
    
endmodule
//
// Verilog Description of module inverter_U563
//

module inverter_U563 (\notGate[491]_keep , \notGate[492] ) /* synthesis syn_module_defined=1 */ ;
    input \notGate[491]_keep ;
    output \notGate[492] ;
    
    wire \notGate[491]_keep  /* synthesis alspreserve=1 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(25[15:22])
    
    LUT4 I1 (.A(\notGate[491]_keep ), .B(\notGate[491]_keep ), .C(\notGate[491]_keep ), 
         .D(\notGate[491]_keep ), .Z(\notGate[492] )) /* synthesis syn_instantiated=1, lut_function=((!D !C !B !A)+(!D !C !B A)+(!D !C B !A)+(!D !C B A)+(!D C !B !A)+(!D C !B A)+(!D C B !A)+(!D C B A)), LSE_LINE_FILE_ID=3, LSE_LCOL=13, LSE_RCOL=44, LSE_LLINE=32, LSE_RLINE=32 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(11[2:53])
    defparam I1.init = 16'b0000000011111111;
    
endmodule
//
// Verilog Description of module inverter_U564
//

module inverter_U564 (\notGate[490]_keep , \notGate[491] ) /* synthesis syn_module_defined=1 */ ;
    input \notGate[490]_keep ;
    output \notGate[491] ;
    
    wire \notGate[490]_keep  /* synthesis alspreserve=1 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(25[15:22])
    
    LUT4 I1 (.A(\notGate[490]_keep ), .B(\notGate[490]_keep ), .C(\notGate[490]_keep ), 
         .D(\notGate[490]_keep ), .Z(\notGate[491] )) /* synthesis syn_instantiated=1, lut_function=((!D !C !B !A)+(!D !C !B A)+(!D !C B !A)+(!D !C B A)+(!D C !B !A)+(!D C !B A)+(!D C B !A)+(!D C B A)), LSE_LINE_FILE_ID=3, LSE_LCOL=13, LSE_RCOL=44, LSE_LLINE=32, LSE_RLINE=32 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(11[2:53])
    defparam I1.init = 16'b0000000011111111;
    
endmodule
//
// Verilog Description of module inverter_U565
//

module inverter_U565 (\notGate[489]_keep , \notGate[490] ) /* synthesis syn_module_defined=1 */ ;
    input \notGate[489]_keep ;
    output \notGate[490] ;
    
    wire \notGate[489]_keep  /* synthesis alspreserve=1 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(25[15:22])
    
    LUT4 I1 (.A(\notGate[489]_keep ), .B(\notGate[489]_keep ), .C(\notGate[489]_keep ), 
         .D(\notGate[489]_keep ), .Z(\notGate[490] )) /* synthesis syn_instantiated=1, lut_function=((!D !C !B !A)+(!D !C !B A)+(!D !C B !A)+(!D !C B A)+(!D C !B !A)+(!D C !B A)+(!D C B !A)+(!D C B A)), LSE_LINE_FILE_ID=3, LSE_LCOL=13, LSE_RCOL=44, LSE_LLINE=32, LSE_RLINE=32 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(11[2:53])
    defparam I1.init = 16'b0000000011111111;
    
endmodule
//
// Verilog Description of module inverter_U566
//

module inverter_U566 (\notGate[47]_keep , \notGate[48] ) /* synthesis syn_module_defined=1 */ ;
    input \notGate[47]_keep ;
    output \notGate[48] ;
    
    wire \notGate[47]_keep  /* synthesis alspreserve=1 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(25[15:22])
    
    LUT4 I1 (.A(\notGate[47]_keep ), .B(\notGate[47]_keep ), .C(\notGate[47]_keep ), 
         .D(\notGate[47]_keep ), .Z(\notGate[48] )) /* synthesis syn_instantiated=1, lut_function=((!D !C !B !A)+(!D !C !B A)+(!D !C B !A)+(!D !C B A)+(!D C !B !A)+(!D C !B A)+(!D C B !A)+(!D C B A)), LSE_LINE_FILE_ID=3, LSE_LCOL=13, LSE_RCOL=44, LSE_LLINE=32, LSE_RLINE=32 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(11[2:53])
    defparam I1.init = 16'b0000000011111111;
    
endmodule
//
// Verilog Description of module inverter_U567
//

module inverter_U567 (\notGate[488]_keep , \notGate[489] ) /* synthesis syn_module_defined=1 */ ;
    input \notGate[488]_keep ;
    output \notGate[489] ;
    
    wire \notGate[488]_keep  /* synthesis alspreserve=1 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(25[15:22])
    
    LUT4 I1 (.A(\notGate[488]_keep ), .B(\notGate[488]_keep ), .C(\notGate[488]_keep ), 
         .D(\notGate[488]_keep ), .Z(\notGate[489] )) /* synthesis syn_instantiated=1, lut_function=((!D !C !B !A)+(!D !C !B A)+(!D !C B !A)+(!D !C B A)+(!D C !B !A)+(!D C !B A)+(!D C B !A)+(!D C B A)), LSE_LINE_FILE_ID=3, LSE_LCOL=13, LSE_RCOL=44, LSE_LLINE=32, LSE_RLINE=32 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(11[2:53])
    defparam I1.init = 16'b0000000011111111;
    
endmodule
//
// Verilog Description of module inverter_U568
//

module inverter_U568 (\notGate[487]_keep , \notGate[488] ) /* synthesis syn_module_defined=1 */ ;
    input \notGate[487]_keep ;
    output \notGate[488] ;
    
    wire \notGate[487]_keep  /* synthesis alspreserve=1 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(25[15:22])
    
    LUT4 I1 (.A(\notGate[487]_keep ), .B(\notGate[487]_keep ), .C(\notGate[487]_keep ), 
         .D(\notGate[487]_keep ), .Z(\notGate[488] )) /* synthesis syn_instantiated=1, lut_function=((!D !C !B !A)+(!D !C !B A)+(!D !C B !A)+(!D !C B A)+(!D C !B !A)+(!D C !B A)+(!D C B !A)+(!D C B A)), LSE_LINE_FILE_ID=3, LSE_LCOL=13, LSE_RCOL=44, LSE_LLINE=32, LSE_RLINE=32 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(11[2:53])
    defparam I1.init = 16'b0000000011111111;
    
endmodule
//
// Verilog Description of module inverter_U569
//

module inverter_U569 (\notGate[486]_keep , \notGate[487] ) /* synthesis syn_module_defined=1 */ ;
    input \notGate[486]_keep ;
    output \notGate[487] ;
    
    wire \notGate[486]_keep  /* synthesis alspreserve=1 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(25[15:22])
    
    LUT4 I1 (.A(\notGate[486]_keep ), .B(\notGate[486]_keep ), .C(\notGate[486]_keep ), 
         .D(\notGate[486]_keep ), .Z(\notGate[487] )) /* synthesis syn_instantiated=1, lut_function=((!D !C !B !A)+(!D !C !B A)+(!D !C B !A)+(!D !C B A)+(!D C !B !A)+(!D C !B A)+(!D C B !A)+(!D C B A)), LSE_LINE_FILE_ID=3, LSE_LCOL=13, LSE_RCOL=44, LSE_LLINE=32, LSE_RLINE=32 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(11[2:53])
    defparam I1.init = 16'b0000000011111111;
    
endmodule
//
// Verilog Description of module inverter_U570
//

module inverter_U570 (\notGate[485]_keep , \notGate[486] ) /* synthesis syn_module_defined=1 */ ;
    input \notGate[485]_keep ;
    output \notGate[486] ;
    
    wire \notGate[485]_keep  /* synthesis alspreserve=1 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(25[15:22])
    
    LUT4 I1 (.A(\notGate[485]_keep ), .B(\notGate[485]_keep ), .C(\notGate[485]_keep ), 
         .D(\notGate[485]_keep ), .Z(\notGate[486] )) /* synthesis syn_instantiated=1, lut_function=((!D !C !B !A)+(!D !C !B A)+(!D !C B !A)+(!D !C B A)+(!D C !B !A)+(!D C !B A)+(!D C B !A)+(!D C B A)), LSE_LINE_FILE_ID=3, LSE_LCOL=13, LSE_RCOL=44, LSE_LLINE=32, LSE_RLINE=32 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(11[2:53])
    defparam I1.init = 16'b0000000011111111;
    
endmodule
//
// Verilog Description of module inverter_U571
//

module inverter_U571 (\notGate[484]_keep , \notGate[485] ) /* synthesis syn_module_defined=1 */ ;
    input \notGate[484]_keep ;
    output \notGate[485] ;
    
    wire \notGate[484]_keep  /* synthesis alspreserve=1 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(25[15:22])
    
    LUT4 I1 (.A(\notGate[484]_keep ), .B(\notGate[484]_keep ), .C(\notGate[484]_keep ), 
         .D(\notGate[484]_keep ), .Z(\notGate[485] )) /* synthesis syn_instantiated=1, lut_function=((!D !C !B !A)+(!D !C !B A)+(!D !C B !A)+(!D !C B A)+(!D C !B !A)+(!D C !B A)+(!D C B !A)+(!D C B A)), LSE_LINE_FILE_ID=3, LSE_LCOL=13, LSE_RCOL=44, LSE_LLINE=32, LSE_RLINE=32 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(11[2:53])
    defparam I1.init = 16'b0000000011111111;
    
endmodule
//
// Verilog Description of module inverter_U572
//

module inverter_U572 (\notGate[483]_keep , \notGate[484] ) /* synthesis syn_module_defined=1 */ ;
    input \notGate[483]_keep ;
    output \notGate[484] ;
    
    wire \notGate[483]_keep  /* synthesis alspreserve=1 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(25[15:22])
    
    LUT4 I1 (.A(\notGate[483]_keep ), .B(\notGate[483]_keep ), .C(\notGate[483]_keep ), 
         .D(\notGate[483]_keep ), .Z(\notGate[484] )) /* synthesis syn_instantiated=1, lut_function=((!D !C !B !A)+(!D !C !B A)+(!D !C B !A)+(!D !C B A)+(!D C !B !A)+(!D C !B A)+(!D C B !A)+(!D C B A)), LSE_LINE_FILE_ID=3, LSE_LCOL=13, LSE_RCOL=44, LSE_LLINE=32, LSE_RLINE=32 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(11[2:53])
    defparam I1.init = 16'b0000000011111111;
    
endmodule
//
// Verilog Description of module inverter_U573
//

module inverter_U573 (\notGate[482]_keep , \notGate[483] ) /* synthesis syn_module_defined=1 */ ;
    input \notGate[482]_keep ;
    output \notGate[483] ;
    
    wire \notGate[482]_keep  /* synthesis alspreserve=1 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(25[15:22])
    
    LUT4 I1 (.A(\notGate[482]_keep ), .B(\notGate[482]_keep ), .C(\notGate[482]_keep ), 
         .D(\notGate[482]_keep ), .Z(\notGate[483] )) /* synthesis syn_instantiated=1, lut_function=((!D !C !B !A)+(!D !C !B A)+(!D !C B !A)+(!D !C B A)+(!D C !B !A)+(!D C !B A)+(!D C B !A)+(!D C B A)), LSE_LINE_FILE_ID=3, LSE_LCOL=13, LSE_RCOL=44, LSE_LLINE=32, LSE_RLINE=32 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(11[2:53])
    defparam I1.init = 16'b0000000011111111;
    
endmodule
//
// Verilog Description of module inverter_U574
//

module inverter_U574 (\notGate[481]_keep , \notGate[482] ) /* synthesis syn_module_defined=1 */ ;
    input \notGate[481]_keep ;
    output \notGate[482] ;
    
    wire \notGate[481]_keep  /* synthesis alspreserve=1 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(25[15:22])
    
    LUT4 I1 (.A(\notGate[481]_keep ), .B(\notGate[481]_keep ), .C(\notGate[481]_keep ), 
         .D(\notGate[481]_keep ), .Z(\notGate[482] )) /* synthesis syn_instantiated=1, lut_function=((!D !C !B !A)+(!D !C !B A)+(!D !C B !A)+(!D !C B A)+(!D C !B !A)+(!D C !B A)+(!D C B !A)+(!D C B A)), LSE_LINE_FILE_ID=3, LSE_LCOL=13, LSE_RCOL=44, LSE_LLINE=32, LSE_RLINE=32 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(11[2:53])
    defparam I1.init = 16'b0000000011111111;
    
endmodule
//
// Verilog Description of module inverter_U575
//

module inverter_U575 (\notGate[480]_keep , \notGate[481] ) /* synthesis syn_module_defined=1 */ ;
    input \notGate[480]_keep ;
    output \notGate[481] ;
    
    wire \notGate[480]_keep  /* synthesis alspreserve=1 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(25[15:22])
    
    LUT4 I1 (.A(\notGate[480]_keep ), .B(\notGate[480]_keep ), .C(\notGate[480]_keep ), 
         .D(\notGate[480]_keep ), .Z(\notGate[481] )) /* synthesis syn_instantiated=1, lut_function=((!D !C !B !A)+(!D !C !B A)+(!D !C B !A)+(!D !C B A)+(!D C !B !A)+(!D C !B A)+(!D C B !A)+(!D C B A)), LSE_LINE_FILE_ID=3, LSE_LCOL=13, LSE_RCOL=44, LSE_LLINE=32, LSE_RLINE=32 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(11[2:53])
    defparam I1.init = 16'b0000000011111111;
    
endmodule
//
// Verilog Description of module inverter_U576
//

module inverter_U576 (\notGate[479]_keep , \notGate[480] ) /* synthesis syn_module_defined=1 */ ;
    input \notGate[479]_keep ;
    output \notGate[480] ;
    
    wire \notGate[479]_keep  /* synthesis alspreserve=1 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(25[15:22])
    
    LUT4 I1 (.A(\notGate[479]_keep ), .B(\notGate[479]_keep ), .C(\notGate[479]_keep ), 
         .D(\notGate[479]_keep ), .Z(\notGate[480] )) /* synthesis syn_instantiated=1, lut_function=((!D !C !B !A)+(!D !C !B A)+(!D !C B !A)+(!D !C B A)+(!D C !B !A)+(!D C !B A)+(!D C B !A)+(!D C B A)), LSE_LINE_FILE_ID=3, LSE_LCOL=13, LSE_RCOL=44, LSE_LLINE=32, LSE_RLINE=32 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(11[2:53])
    defparam I1.init = 16'b0000000011111111;
    
endmodule
//
// Verilog Description of module inverter_U577
//

module inverter_U577 (\notGate[46]_keep , \notGate[47] ) /* synthesis syn_module_defined=1 */ ;
    input \notGate[46]_keep ;
    output \notGate[47] ;
    
    wire \notGate[46]_keep  /* synthesis alspreserve=1 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(25[15:22])
    
    LUT4 I1 (.A(\notGate[46]_keep ), .B(\notGate[46]_keep ), .C(\notGate[46]_keep ), 
         .D(\notGate[46]_keep ), .Z(\notGate[47] )) /* synthesis syn_instantiated=1, lut_function=((!D !C !B !A)+(!D !C !B A)+(!D !C B !A)+(!D !C B A)+(!D C !B !A)+(!D C !B A)+(!D C B !A)+(!D C B A)), LSE_LINE_FILE_ID=3, LSE_LCOL=13, LSE_RCOL=44, LSE_LLINE=32, LSE_RLINE=32 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(11[2:53])
    defparam I1.init = 16'b0000000011111111;
    
endmodule
//
// Verilog Description of module inverter_U578
//

module inverter_U578 (\notGate[478]_keep , \notGate[479] ) /* synthesis syn_module_defined=1 */ ;
    input \notGate[478]_keep ;
    output \notGate[479] ;
    
    wire \notGate[478]_keep  /* synthesis alspreserve=1 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(25[15:22])
    
    LUT4 I1 (.A(\notGate[478]_keep ), .B(\notGate[478]_keep ), .C(\notGate[478]_keep ), 
         .D(\notGate[478]_keep ), .Z(\notGate[479] )) /* synthesis syn_instantiated=1, lut_function=((!D !C !B !A)+(!D !C !B A)+(!D !C B !A)+(!D !C B A)+(!D C !B !A)+(!D C !B A)+(!D C B !A)+(!D C B A)), LSE_LINE_FILE_ID=3, LSE_LCOL=13, LSE_RCOL=44, LSE_LLINE=32, LSE_RLINE=32 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(11[2:53])
    defparam I1.init = 16'b0000000011111111;
    
endmodule
//
// Verilog Description of module inverter_U579
//

module inverter_U579 (\notGate[477]_keep , \notGate[478] ) /* synthesis syn_module_defined=1 */ ;
    input \notGate[477]_keep ;
    output \notGate[478] ;
    
    wire \notGate[477]_keep  /* synthesis alspreserve=1 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(25[15:22])
    
    LUT4 I1 (.A(\notGate[477]_keep ), .B(\notGate[477]_keep ), .C(\notGate[477]_keep ), 
         .D(\notGate[477]_keep ), .Z(\notGate[478] )) /* synthesis syn_instantiated=1, lut_function=((!D !C !B !A)+(!D !C !B A)+(!D !C B !A)+(!D !C B A)+(!D C !B !A)+(!D C !B A)+(!D C B !A)+(!D C B A)), LSE_LINE_FILE_ID=3, LSE_LCOL=13, LSE_RCOL=44, LSE_LLINE=32, LSE_RLINE=32 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(11[2:53])
    defparam I1.init = 16'b0000000011111111;
    
endmodule
//
// Verilog Description of module inverter_U580
//

module inverter_U580 (\notGate[476]_keep , \notGate[477] ) /* synthesis syn_module_defined=1 */ ;
    input \notGate[476]_keep ;
    output \notGate[477] ;
    
    wire \notGate[476]_keep  /* synthesis alspreserve=1 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(25[15:22])
    
    LUT4 I1 (.A(\notGate[476]_keep ), .B(\notGate[476]_keep ), .C(\notGate[476]_keep ), 
         .D(\notGate[476]_keep ), .Z(\notGate[477] )) /* synthesis syn_instantiated=1, lut_function=((!D !C !B !A)+(!D !C !B A)+(!D !C B !A)+(!D !C B A)+(!D C !B !A)+(!D C !B A)+(!D C B !A)+(!D C B A)), LSE_LINE_FILE_ID=3, LSE_LCOL=13, LSE_RCOL=44, LSE_LLINE=32, LSE_RLINE=32 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(11[2:53])
    defparam I1.init = 16'b0000000011111111;
    
endmodule
//
// Verilog Description of module inverter_U581
//

module inverter_U581 (\notGate[475]_keep , \notGate[476] ) /* synthesis syn_module_defined=1 */ ;
    input \notGate[475]_keep ;
    output \notGate[476] ;
    
    wire \notGate[475]_keep  /* synthesis alspreserve=1 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(25[15:22])
    
    LUT4 I1 (.A(\notGate[475]_keep ), .B(\notGate[475]_keep ), .C(\notGate[475]_keep ), 
         .D(\notGate[475]_keep ), .Z(\notGate[476] )) /* synthesis syn_instantiated=1, lut_function=((!D !C !B !A)+(!D !C !B A)+(!D !C B !A)+(!D !C B A)+(!D C !B !A)+(!D C !B A)+(!D C B !A)+(!D C B A)), LSE_LINE_FILE_ID=3, LSE_LCOL=13, LSE_RCOL=44, LSE_LLINE=32, LSE_RLINE=32 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(11[2:53])
    defparam I1.init = 16'b0000000011111111;
    
endmodule
//
// Verilog Description of module inverter_U582
//

module inverter_U582 (\notGate[474]_keep , \notGate[475] ) /* synthesis syn_module_defined=1 */ ;
    input \notGate[474]_keep ;
    output \notGate[475] ;
    
    wire \notGate[474]_keep  /* synthesis alspreserve=1 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(25[15:22])
    
    LUT4 I1 (.A(\notGate[474]_keep ), .B(\notGate[474]_keep ), .C(\notGate[474]_keep ), 
         .D(\notGate[474]_keep ), .Z(\notGate[475] )) /* synthesis syn_instantiated=1, lut_function=((!D !C !B !A)+(!D !C !B A)+(!D !C B !A)+(!D !C B A)+(!D C !B !A)+(!D C !B A)+(!D C B !A)+(!D C B A)), LSE_LINE_FILE_ID=3, LSE_LCOL=13, LSE_RCOL=44, LSE_LLINE=32, LSE_RLINE=32 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(11[2:53])
    defparam I1.init = 16'b0000000011111111;
    
endmodule
//
// Verilog Description of module inverter_U583
//

module inverter_U583 (\notGate[473]_keep , \notGate[474] ) /* synthesis syn_module_defined=1 */ ;
    input \notGate[473]_keep ;
    output \notGate[474] ;
    
    wire \notGate[473]_keep  /* synthesis alspreserve=1 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(25[15:22])
    
    LUT4 I1 (.A(\notGate[473]_keep ), .B(\notGate[473]_keep ), .C(\notGate[473]_keep ), 
         .D(\notGate[473]_keep ), .Z(\notGate[474] )) /* synthesis syn_instantiated=1, lut_function=((!D !C !B !A)+(!D !C !B A)+(!D !C B !A)+(!D !C B A)+(!D C !B !A)+(!D C !B A)+(!D C B !A)+(!D C B A)), LSE_LINE_FILE_ID=3, LSE_LCOL=13, LSE_RCOL=44, LSE_LLINE=32, LSE_RLINE=32 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(11[2:53])
    defparam I1.init = 16'b0000000011111111;
    
endmodule
//
// Verilog Description of module inverter_U584
//

module inverter_U584 (\notGate[472]_keep , \notGate[473] ) /* synthesis syn_module_defined=1 */ ;
    input \notGate[472]_keep ;
    output \notGate[473] ;
    
    wire \notGate[472]_keep  /* synthesis alspreserve=1 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(25[15:22])
    
    LUT4 I1 (.A(\notGate[472]_keep ), .B(\notGate[472]_keep ), .C(\notGate[472]_keep ), 
         .D(\notGate[472]_keep ), .Z(\notGate[473] )) /* synthesis syn_instantiated=1, lut_function=((!D !C !B !A)+(!D !C !B A)+(!D !C B !A)+(!D !C B A)+(!D C !B !A)+(!D C !B A)+(!D C B !A)+(!D C B A)), LSE_LINE_FILE_ID=3, LSE_LCOL=13, LSE_RCOL=44, LSE_LLINE=32, LSE_RLINE=32 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(11[2:53])
    defparam I1.init = 16'b0000000011111111;
    
endmodule
//
// Verilog Description of module inverter_U585
//

module inverter_U585 (\notGate[471]_keep , \notGate[472] ) /* synthesis syn_module_defined=1 */ ;
    input \notGate[471]_keep ;
    output \notGate[472] ;
    
    wire \notGate[471]_keep  /* synthesis alspreserve=1 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(25[15:22])
    
    LUT4 I1 (.A(\notGate[471]_keep ), .B(\notGate[471]_keep ), .C(\notGate[471]_keep ), 
         .D(\notGate[471]_keep ), .Z(\notGate[472] )) /* synthesis syn_instantiated=1, lut_function=((!D !C !B !A)+(!D !C !B A)+(!D !C B !A)+(!D !C B A)+(!D C !B !A)+(!D C !B A)+(!D C B !A)+(!D C B A)), LSE_LINE_FILE_ID=3, LSE_LCOL=13, LSE_RCOL=44, LSE_LLINE=32, LSE_RLINE=32 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(11[2:53])
    defparam I1.init = 16'b0000000011111111;
    
endmodule
//
// Verilog Description of module inverter_U586
//

module inverter_U586 (\notGate[470]_keep , \notGate[471] ) /* synthesis syn_module_defined=1 */ ;
    input \notGate[470]_keep ;
    output \notGate[471] ;
    
    wire \notGate[470]_keep  /* synthesis alspreserve=1 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(25[15:22])
    
    LUT4 I1 (.A(\notGate[470]_keep ), .B(\notGate[470]_keep ), .C(\notGate[470]_keep ), 
         .D(\notGate[470]_keep ), .Z(\notGate[471] )) /* synthesis syn_instantiated=1, lut_function=((!D !C !B !A)+(!D !C !B A)+(!D !C B !A)+(!D !C B A)+(!D C !B !A)+(!D C !B A)+(!D C B !A)+(!D C B A)), LSE_LINE_FILE_ID=3, LSE_LCOL=13, LSE_RCOL=44, LSE_LLINE=32, LSE_RLINE=32 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(11[2:53])
    defparam I1.init = 16'b0000000011111111;
    
endmodule
//
// Verilog Description of module inverter_U587
//

module inverter_U587 (\notGate[469]_keep , \notGate[470] ) /* synthesis syn_module_defined=1 */ ;
    input \notGate[469]_keep ;
    output \notGate[470] ;
    
    wire \notGate[469]_keep  /* synthesis alspreserve=1 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(25[15:22])
    
    LUT4 I1 (.A(\notGate[469]_keep ), .B(\notGate[469]_keep ), .C(\notGate[469]_keep ), 
         .D(\notGate[469]_keep ), .Z(\notGate[470] )) /* synthesis syn_instantiated=1, lut_function=((!D !C !B !A)+(!D !C !B A)+(!D !C B !A)+(!D !C B A)+(!D C !B !A)+(!D C !B A)+(!D C B !A)+(!D C B A)), LSE_LINE_FILE_ID=3, LSE_LCOL=13, LSE_RCOL=44, LSE_LLINE=32, LSE_RLINE=32 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(11[2:53])
    defparam I1.init = 16'b0000000011111111;
    
endmodule
//
// Verilog Description of module inverter_U588
//

module inverter_U588 (\notGate[45]_keep , \notGate[46] ) /* synthesis syn_module_defined=1 */ ;
    input \notGate[45]_keep ;
    output \notGate[46] ;
    
    wire \notGate[45]_keep  /* synthesis alspreserve=1 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(25[15:22])
    
    LUT4 I1 (.A(\notGate[45]_keep ), .B(\notGate[45]_keep ), .C(\notGate[45]_keep ), 
         .D(\notGate[45]_keep ), .Z(\notGate[46] )) /* synthesis syn_instantiated=1, lut_function=((!D !C !B !A)+(!D !C !B A)+(!D !C B !A)+(!D !C B A)+(!D C !B !A)+(!D C !B A)+(!D C B !A)+(!D C B A)), LSE_LINE_FILE_ID=3, LSE_LCOL=13, LSE_RCOL=44, LSE_LLINE=32, LSE_RLINE=32 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(11[2:53])
    defparam I1.init = 16'b0000000011111111;
    
endmodule
//
// Verilog Description of module inverter_U589
//

module inverter_U589 (\notGate[468]_keep , \notGate[469] ) /* synthesis syn_module_defined=1 */ ;
    input \notGate[468]_keep ;
    output \notGate[469] ;
    
    wire \notGate[468]_keep  /* synthesis alspreserve=1 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(25[15:22])
    
    LUT4 I1 (.A(\notGate[468]_keep ), .B(\notGate[468]_keep ), .C(\notGate[468]_keep ), 
         .D(\notGate[468]_keep ), .Z(\notGate[469] )) /* synthesis syn_instantiated=1, lut_function=((!D !C !B !A)+(!D !C !B A)+(!D !C B !A)+(!D !C B A)+(!D C !B !A)+(!D C !B A)+(!D C B !A)+(!D C B A)), LSE_LINE_FILE_ID=3, LSE_LCOL=13, LSE_RCOL=44, LSE_LLINE=32, LSE_RLINE=32 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(11[2:53])
    defparam I1.init = 16'b0000000011111111;
    
endmodule
//
// Verilog Description of module inverter_U590
//

module inverter_U590 (\notGate[467]_keep , \notGate[468] ) /* synthesis syn_module_defined=1 */ ;
    input \notGate[467]_keep ;
    output \notGate[468] ;
    
    wire \notGate[467]_keep  /* synthesis alspreserve=1 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(25[15:22])
    
    LUT4 I1 (.A(\notGate[467]_keep ), .B(\notGate[467]_keep ), .C(\notGate[467]_keep ), 
         .D(\notGate[467]_keep ), .Z(\notGate[468] )) /* synthesis syn_instantiated=1, lut_function=((!D !C !B !A)+(!D !C !B A)+(!D !C B !A)+(!D !C B A)+(!D C !B !A)+(!D C !B A)+(!D C B !A)+(!D C B A)), LSE_LINE_FILE_ID=3, LSE_LCOL=13, LSE_RCOL=44, LSE_LLINE=32, LSE_RLINE=32 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(11[2:53])
    defparam I1.init = 16'b0000000011111111;
    
endmodule
//
// Verilog Description of module inverter_U591
//

module inverter_U591 (\notGate[466]_keep , \notGate[467] ) /* synthesis syn_module_defined=1 */ ;
    input \notGate[466]_keep ;
    output \notGate[467] ;
    
    wire \notGate[466]_keep  /* synthesis alspreserve=1 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(25[15:22])
    
    LUT4 I1 (.A(\notGate[466]_keep ), .B(\notGate[466]_keep ), .C(\notGate[466]_keep ), 
         .D(\notGate[466]_keep ), .Z(\notGate[467] )) /* synthesis syn_instantiated=1, lut_function=((!D !C !B !A)+(!D !C !B A)+(!D !C B !A)+(!D !C B A)+(!D C !B !A)+(!D C !B A)+(!D C B !A)+(!D C B A)), LSE_LINE_FILE_ID=3, LSE_LCOL=13, LSE_RCOL=44, LSE_LLINE=32, LSE_RLINE=32 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(11[2:53])
    defparam I1.init = 16'b0000000011111111;
    
endmodule
//
// Verilog Description of module inverter_U592
//

module inverter_U592 (\notGate[465]_keep , \notGate[466] ) /* synthesis syn_module_defined=1 */ ;
    input \notGate[465]_keep ;
    output \notGate[466] ;
    
    wire \notGate[465]_keep  /* synthesis alspreserve=1 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(25[15:22])
    
    LUT4 I1 (.A(\notGate[465]_keep ), .B(\notGate[465]_keep ), .C(\notGate[465]_keep ), 
         .D(\notGate[465]_keep ), .Z(\notGate[466] )) /* synthesis syn_instantiated=1, lut_function=((!D !C !B !A)+(!D !C !B A)+(!D !C B !A)+(!D !C B A)+(!D C !B !A)+(!D C !B A)+(!D C B !A)+(!D C B A)), LSE_LINE_FILE_ID=3, LSE_LCOL=13, LSE_RCOL=44, LSE_LLINE=32, LSE_RLINE=32 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(11[2:53])
    defparam I1.init = 16'b0000000011111111;
    
endmodule
//
// Verilog Description of module inverter_U593
//

module inverter_U593 (\notGate[464]_keep , \notGate[465] ) /* synthesis syn_module_defined=1 */ ;
    input \notGate[464]_keep ;
    output \notGate[465] ;
    
    wire \notGate[464]_keep  /* synthesis alspreserve=1 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(25[15:22])
    
    LUT4 I1 (.A(\notGate[464]_keep ), .B(\notGate[464]_keep ), .C(\notGate[464]_keep ), 
         .D(\notGate[464]_keep ), .Z(\notGate[465] )) /* synthesis syn_instantiated=1, lut_function=((!D !C !B !A)+(!D !C !B A)+(!D !C B !A)+(!D !C B A)+(!D C !B !A)+(!D C !B A)+(!D C B !A)+(!D C B A)), LSE_LINE_FILE_ID=3, LSE_LCOL=13, LSE_RCOL=44, LSE_LLINE=32, LSE_RLINE=32 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(11[2:53])
    defparam I1.init = 16'b0000000011111111;
    
endmodule
//
// Verilog Description of module inverter_U594
//

module inverter_U594 (\notGate[463]_keep , \notGate[464] ) /* synthesis syn_module_defined=1 */ ;
    input \notGate[463]_keep ;
    output \notGate[464] ;
    
    wire \notGate[463]_keep  /* synthesis alspreserve=1 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(25[15:22])
    
    LUT4 I1 (.A(\notGate[463]_keep ), .B(\notGate[463]_keep ), .C(\notGate[463]_keep ), 
         .D(\notGate[463]_keep ), .Z(\notGate[464] )) /* synthesis syn_instantiated=1, lut_function=((!D !C !B !A)+(!D !C !B A)+(!D !C B !A)+(!D !C B A)+(!D C !B !A)+(!D C !B A)+(!D C B !A)+(!D C B A)), LSE_LINE_FILE_ID=3, LSE_LCOL=13, LSE_RCOL=44, LSE_LLINE=32, LSE_RLINE=32 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(11[2:53])
    defparam I1.init = 16'b0000000011111111;
    
endmodule
//
// Verilog Description of module inverter_U595
//

module inverter_U595 (\notGate[462]_keep , \notGate[463] ) /* synthesis syn_module_defined=1 */ ;
    input \notGate[462]_keep ;
    output \notGate[463] ;
    
    wire \notGate[462]_keep  /* synthesis alspreserve=1 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(25[15:22])
    
    LUT4 I1 (.A(\notGate[462]_keep ), .B(\notGate[462]_keep ), .C(\notGate[462]_keep ), 
         .D(\notGate[462]_keep ), .Z(\notGate[463] )) /* synthesis syn_instantiated=1, lut_function=((!D !C !B !A)+(!D !C !B A)+(!D !C B !A)+(!D !C B A)+(!D C !B !A)+(!D C !B A)+(!D C B !A)+(!D C B A)), LSE_LINE_FILE_ID=3, LSE_LCOL=13, LSE_RCOL=44, LSE_LLINE=32, LSE_RLINE=32 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(11[2:53])
    defparam I1.init = 16'b0000000011111111;
    
endmodule
//
// Verilog Description of module inverter_U596
//

module inverter_U596 (\notGate[461]_keep , \notGate[462] ) /* synthesis syn_module_defined=1 */ ;
    input \notGate[461]_keep ;
    output \notGate[462] ;
    
    wire \notGate[461]_keep  /* synthesis alspreserve=1 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(25[15:22])
    
    LUT4 I1 (.A(\notGate[461]_keep ), .B(\notGate[461]_keep ), .C(\notGate[461]_keep ), 
         .D(\notGate[461]_keep ), .Z(\notGate[462] )) /* synthesis syn_instantiated=1, lut_function=((!D !C !B !A)+(!D !C !B A)+(!D !C B !A)+(!D !C B A)+(!D C !B !A)+(!D C !B A)+(!D C B !A)+(!D C B A)), LSE_LINE_FILE_ID=3, LSE_LCOL=13, LSE_RCOL=44, LSE_LLINE=32, LSE_RLINE=32 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(11[2:53])
    defparam I1.init = 16'b0000000011111111;
    
endmodule
//
// Verilog Description of module inverter_U597
//

module inverter_U597 (\notGate[460]_keep , \notGate[461] ) /* synthesis syn_module_defined=1 */ ;
    input \notGate[460]_keep ;
    output \notGate[461] ;
    
    wire \notGate[460]_keep  /* synthesis alspreserve=1 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(25[15:22])
    
    LUT4 I1 (.A(\notGate[460]_keep ), .B(\notGate[460]_keep ), .C(\notGate[460]_keep ), 
         .D(\notGate[460]_keep ), .Z(\notGate[461] )) /* synthesis syn_instantiated=1, lut_function=((!D !C !B !A)+(!D !C !B A)+(!D !C B !A)+(!D !C B A)+(!D C !B !A)+(!D C !B A)+(!D C B !A)+(!D C B A)), LSE_LINE_FILE_ID=3, LSE_LCOL=13, LSE_RCOL=44, LSE_LLINE=32, LSE_RLINE=32 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(11[2:53])
    defparam I1.init = 16'b0000000011111111;
    
endmodule
//
// Verilog Description of module inverter_U598
//

module inverter_U598 (\notGate[459]_keep , \notGate[460] ) /* synthesis syn_module_defined=1 */ ;
    input \notGate[459]_keep ;
    output \notGate[460] ;
    
    wire \notGate[459]_keep  /* synthesis alspreserve=1 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(25[15:22])
    
    LUT4 I1 (.A(\notGate[459]_keep ), .B(\notGate[459]_keep ), .C(\notGate[459]_keep ), 
         .D(\notGate[459]_keep ), .Z(\notGate[460] )) /* synthesis syn_instantiated=1, lut_function=((!D !C !B !A)+(!D !C !B A)+(!D !C B !A)+(!D !C B A)+(!D C !B !A)+(!D C !B A)+(!D C B !A)+(!D C B A)), LSE_LINE_FILE_ID=3, LSE_LCOL=13, LSE_RCOL=44, LSE_LLINE=32, LSE_RLINE=32 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(11[2:53])
    defparam I1.init = 16'b0000000011111111;
    
endmodule
//
// Verilog Description of module inverter_U599
//

module inverter_U599 (\notGate[44]_keep , \notGate[45] ) /* synthesis syn_module_defined=1 */ ;
    input \notGate[44]_keep ;
    output \notGate[45] ;
    
    wire \notGate[44]_keep  /* synthesis alspreserve=1 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(25[15:22])
    
    LUT4 I1 (.A(\notGate[44]_keep ), .B(\notGate[44]_keep ), .C(\notGate[44]_keep ), 
         .D(\notGate[44]_keep ), .Z(\notGate[45] )) /* synthesis syn_instantiated=1, lut_function=((!D !C !B !A)+(!D !C !B A)+(!D !C B !A)+(!D !C B A)+(!D C !B !A)+(!D C !B A)+(!D C B !A)+(!D C B A)), LSE_LINE_FILE_ID=3, LSE_LCOL=13, LSE_RCOL=44, LSE_LLINE=32, LSE_RLINE=32 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(11[2:53])
    defparam I1.init = 16'b0000000011111111;
    
endmodule
//
// Verilog Description of module inverter_U600
//

module inverter_U600 (\notGate[458]_keep , \notGate[459] ) /* synthesis syn_module_defined=1 */ ;
    input \notGate[458]_keep ;
    output \notGate[459] ;
    
    wire \notGate[458]_keep  /* synthesis alspreserve=1 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(25[15:22])
    
    LUT4 I1 (.A(\notGate[458]_keep ), .B(\notGate[458]_keep ), .C(\notGate[458]_keep ), 
         .D(\notGate[458]_keep ), .Z(\notGate[459] )) /* synthesis syn_instantiated=1, lut_function=((!D !C !B !A)+(!D !C !B A)+(!D !C B !A)+(!D !C B A)+(!D C !B !A)+(!D C !B A)+(!D C B !A)+(!D C B A)), LSE_LINE_FILE_ID=3, LSE_LCOL=13, LSE_RCOL=44, LSE_LLINE=32, LSE_RLINE=32 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(11[2:53])
    defparam I1.init = 16'b0000000011111111;
    
endmodule
//
// Verilog Description of module inverter_U601
//

module inverter_U601 (\notGate[457]_keep , \notGate[458] ) /* synthesis syn_module_defined=1 */ ;
    input \notGate[457]_keep ;
    output \notGate[458] ;
    
    wire \notGate[457]_keep  /* synthesis alspreserve=1 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(25[15:22])
    
    LUT4 I1 (.A(\notGate[457]_keep ), .B(\notGate[457]_keep ), .C(\notGate[457]_keep ), 
         .D(\notGate[457]_keep ), .Z(\notGate[458] )) /* synthesis syn_instantiated=1, lut_function=((!D !C !B !A)+(!D !C !B A)+(!D !C B !A)+(!D !C B A)+(!D C !B !A)+(!D C !B A)+(!D C B !A)+(!D C B A)), LSE_LINE_FILE_ID=3, LSE_LCOL=13, LSE_RCOL=44, LSE_LLINE=32, LSE_RLINE=32 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(11[2:53])
    defparam I1.init = 16'b0000000011111111;
    
endmodule
//
// Verilog Description of module inverter_U602
//

module inverter_U602 (\notGate[456]_keep , \notGate[457] ) /* synthesis syn_module_defined=1 */ ;
    input \notGate[456]_keep ;
    output \notGate[457] ;
    
    wire \notGate[456]_keep  /* synthesis alspreserve=1 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(25[15:22])
    
    LUT4 I1 (.A(\notGate[456]_keep ), .B(\notGate[456]_keep ), .C(\notGate[456]_keep ), 
         .D(\notGate[456]_keep ), .Z(\notGate[457] )) /* synthesis syn_instantiated=1, lut_function=((!D !C !B !A)+(!D !C !B A)+(!D !C B !A)+(!D !C B A)+(!D C !B !A)+(!D C !B A)+(!D C B !A)+(!D C B A)), LSE_LINE_FILE_ID=3, LSE_LCOL=13, LSE_RCOL=44, LSE_LLINE=32, LSE_RLINE=32 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(11[2:53])
    defparam I1.init = 16'b0000000011111111;
    
endmodule
//
// Verilog Description of module inverter_U603
//

module inverter_U603 (\notGate[455]_keep , \notGate[456] ) /* synthesis syn_module_defined=1 */ ;
    input \notGate[455]_keep ;
    output \notGate[456] ;
    
    wire \notGate[455]_keep  /* synthesis alspreserve=1 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(25[15:22])
    
    LUT4 I1 (.A(\notGate[455]_keep ), .B(\notGate[455]_keep ), .C(\notGate[455]_keep ), 
         .D(\notGate[455]_keep ), .Z(\notGate[456] )) /* synthesis syn_instantiated=1, lut_function=((!D !C !B !A)+(!D !C !B A)+(!D !C B !A)+(!D !C B A)+(!D C !B !A)+(!D C !B A)+(!D C B !A)+(!D C B A)), LSE_LINE_FILE_ID=3, LSE_LCOL=13, LSE_RCOL=44, LSE_LLINE=32, LSE_RLINE=32 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(11[2:53])
    defparam I1.init = 16'b0000000011111111;
    
endmodule
//
// Verilog Description of module inverter_U604
//

module inverter_U604 (\notGate[454]_keep , \notGate[455] ) /* synthesis syn_module_defined=1 */ ;
    input \notGate[454]_keep ;
    output \notGate[455] ;
    
    wire \notGate[454]_keep  /* synthesis alspreserve=1 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(25[15:22])
    
    LUT4 I1 (.A(\notGate[454]_keep ), .B(\notGate[454]_keep ), .C(\notGate[454]_keep ), 
         .D(\notGate[454]_keep ), .Z(\notGate[455] )) /* synthesis syn_instantiated=1, lut_function=((!D !C !B !A)+(!D !C !B A)+(!D !C B !A)+(!D !C B A)+(!D C !B !A)+(!D C !B A)+(!D C B !A)+(!D C B A)), LSE_LINE_FILE_ID=3, LSE_LCOL=13, LSE_RCOL=44, LSE_LLINE=32, LSE_RLINE=32 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(11[2:53])
    defparam I1.init = 16'b0000000011111111;
    
endmodule
//
// Verilog Description of module inverter_U605
//

module inverter_U605 (\notGate[453]_keep , \notGate[454] ) /* synthesis syn_module_defined=1 */ ;
    input \notGate[453]_keep ;
    output \notGate[454] ;
    
    wire \notGate[453]_keep  /* synthesis alspreserve=1 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(25[15:22])
    
    LUT4 I1 (.A(\notGate[453]_keep ), .B(\notGate[453]_keep ), .C(\notGate[453]_keep ), 
         .D(\notGate[453]_keep ), .Z(\notGate[454] )) /* synthesis syn_instantiated=1, lut_function=((!D !C !B !A)+(!D !C !B A)+(!D !C B !A)+(!D !C B A)+(!D C !B !A)+(!D C !B A)+(!D C B !A)+(!D C B A)), LSE_LINE_FILE_ID=3, LSE_LCOL=13, LSE_RCOL=44, LSE_LLINE=32, LSE_RLINE=32 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(11[2:53])
    defparam I1.init = 16'b0000000011111111;
    
endmodule
//
// Verilog Description of module inverter_U606
//

module inverter_U606 (\notGate[452]_keep , \notGate[453] ) /* synthesis syn_module_defined=1 */ ;
    input \notGate[452]_keep ;
    output \notGate[453] ;
    
    wire \notGate[452]_keep  /* synthesis alspreserve=1 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(25[15:22])
    
    LUT4 I1 (.A(\notGate[452]_keep ), .B(\notGate[452]_keep ), .C(\notGate[452]_keep ), 
         .D(\notGate[452]_keep ), .Z(\notGate[453] )) /* synthesis syn_instantiated=1, lut_function=((!D !C !B !A)+(!D !C !B A)+(!D !C B !A)+(!D !C B A)+(!D C !B !A)+(!D C !B A)+(!D C B !A)+(!D C B A)), LSE_LINE_FILE_ID=3, LSE_LCOL=13, LSE_RCOL=44, LSE_LLINE=32, LSE_RLINE=32 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(11[2:53])
    defparam I1.init = 16'b0000000011111111;
    
endmodule
//
// Verilog Description of module inverter_U607
//

module inverter_U607 (\notGate[451]_keep , \notGate[452] ) /* synthesis syn_module_defined=1 */ ;
    input \notGate[451]_keep ;
    output \notGate[452] ;
    
    wire \notGate[451]_keep  /* synthesis alspreserve=1 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(25[15:22])
    
    LUT4 I1 (.A(\notGate[451]_keep ), .B(\notGate[451]_keep ), .C(\notGate[451]_keep ), 
         .D(\notGate[451]_keep ), .Z(\notGate[452] )) /* synthesis syn_instantiated=1, lut_function=((!D !C !B !A)+(!D !C !B A)+(!D !C B !A)+(!D !C B A)+(!D C !B !A)+(!D C !B A)+(!D C B !A)+(!D C B A)), LSE_LINE_FILE_ID=3, LSE_LCOL=13, LSE_RCOL=44, LSE_LLINE=32, LSE_RLINE=32 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(11[2:53])
    defparam I1.init = 16'b0000000011111111;
    
endmodule
//
// Verilog Description of module inverter_U608
//

module inverter_U608 (\notGate[450]_keep , \notGate[451] ) /* synthesis syn_module_defined=1 */ ;
    input \notGate[450]_keep ;
    output \notGate[451] ;
    
    wire \notGate[450]_keep  /* synthesis alspreserve=1 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(25[15:22])
    
    LUT4 I1 (.A(\notGate[450]_keep ), .B(\notGate[450]_keep ), .C(\notGate[450]_keep ), 
         .D(\notGate[450]_keep ), .Z(\notGate[451] )) /* synthesis syn_instantiated=1, lut_function=((!D !C !B !A)+(!D !C !B A)+(!D !C B !A)+(!D !C B A)+(!D C !B !A)+(!D C !B A)+(!D C B !A)+(!D C B A)), LSE_LINE_FILE_ID=3, LSE_LCOL=13, LSE_RCOL=44, LSE_LLINE=32, LSE_RLINE=32 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(11[2:53])
    defparam I1.init = 16'b0000000011111111;
    
endmodule
//
// Verilog Description of module inverter_U609
//

module inverter_U609 (\notGate[449]_keep , \notGate[450] ) /* synthesis syn_module_defined=1 */ ;
    input \notGate[449]_keep ;
    output \notGate[450] ;
    
    wire \notGate[449]_keep  /* synthesis alspreserve=1 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(25[15:22])
    
    LUT4 I1 (.A(\notGate[449]_keep ), .B(\notGate[449]_keep ), .C(\notGate[449]_keep ), 
         .D(\notGate[449]_keep ), .Z(\notGate[450] )) /* synthesis syn_instantiated=1, lut_function=((!D !C !B !A)+(!D !C !B A)+(!D !C B !A)+(!D !C B A)+(!D C !B !A)+(!D C !B A)+(!D C B !A)+(!D C B A)), LSE_LINE_FILE_ID=3, LSE_LCOL=13, LSE_RCOL=44, LSE_LLINE=32, LSE_RLINE=32 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(11[2:53])
    defparam I1.init = 16'b0000000011111111;
    
endmodule
//
// Verilog Description of module inverter_U610
//

module inverter_U610 (\notGate[43]_keep , \notGate[44] ) /* synthesis syn_module_defined=1 */ ;
    input \notGate[43]_keep ;
    output \notGate[44] ;
    
    wire \notGate[43]_keep  /* synthesis alspreserve=1 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(25[15:22])
    
    LUT4 I1 (.A(\notGate[43]_keep ), .B(\notGate[43]_keep ), .C(\notGate[43]_keep ), 
         .D(\notGate[43]_keep ), .Z(\notGate[44] )) /* synthesis syn_instantiated=1, lut_function=((!D !C !B !A)+(!D !C !B A)+(!D !C B !A)+(!D !C B A)+(!D C !B !A)+(!D C !B A)+(!D C B !A)+(!D C B A)), LSE_LINE_FILE_ID=3, LSE_LCOL=13, LSE_RCOL=44, LSE_LLINE=32, LSE_RLINE=32 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(11[2:53])
    defparam I1.init = 16'b0000000011111111;
    
endmodule
//
// Verilog Description of module inverter_U611
//

module inverter_U611 (\notGate[448]_keep , \notGate[449] ) /* synthesis syn_module_defined=1 */ ;
    input \notGate[448]_keep ;
    output \notGate[449] ;
    
    wire \notGate[448]_keep  /* synthesis alspreserve=1 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(25[15:22])
    
    LUT4 I1 (.A(\notGate[448]_keep ), .B(\notGate[448]_keep ), .C(\notGate[448]_keep ), 
         .D(\notGate[448]_keep ), .Z(\notGate[449] )) /* synthesis syn_instantiated=1, lut_function=((!D !C !B !A)+(!D !C !B A)+(!D !C B !A)+(!D !C B A)+(!D C !B !A)+(!D C !B A)+(!D C B !A)+(!D C B A)), LSE_LINE_FILE_ID=3, LSE_LCOL=13, LSE_RCOL=44, LSE_LLINE=32, LSE_RLINE=32 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(11[2:53])
    defparam I1.init = 16'b0000000011111111;
    
endmodule
//
// Verilog Description of module inverter_U612
//

module inverter_U612 (\notGate[447]_keep , \notGate[448] ) /* synthesis syn_module_defined=1 */ ;
    input \notGate[447]_keep ;
    output \notGate[448] ;
    
    wire \notGate[447]_keep  /* synthesis alspreserve=1 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(25[15:22])
    
    LUT4 I1 (.A(\notGate[447]_keep ), .B(\notGate[447]_keep ), .C(\notGate[447]_keep ), 
         .D(\notGate[447]_keep ), .Z(\notGate[448] )) /* synthesis syn_instantiated=1, lut_function=((!D !C !B !A)+(!D !C !B A)+(!D !C B !A)+(!D !C B A)+(!D C !B !A)+(!D C !B A)+(!D C B !A)+(!D C B A)), LSE_LINE_FILE_ID=3, LSE_LCOL=13, LSE_RCOL=44, LSE_LLINE=32, LSE_RLINE=32 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(11[2:53])
    defparam I1.init = 16'b0000000011111111;
    
endmodule
//
// Verilog Description of module inverter_U613
//

module inverter_U613 (\notGate[446]_keep , \notGate[447] ) /* synthesis syn_module_defined=1 */ ;
    input \notGate[446]_keep ;
    output \notGate[447] ;
    
    wire \notGate[446]_keep  /* synthesis alspreserve=1 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(25[15:22])
    
    LUT4 I1 (.A(\notGate[446]_keep ), .B(\notGate[446]_keep ), .C(\notGate[446]_keep ), 
         .D(\notGate[446]_keep ), .Z(\notGate[447] )) /* synthesis syn_instantiated=1, lut_function=((!D !C !B !A)+(!D !C !B A)+(!D !C B !A)+(!D !C B A)+(!D C !B !A)+(!D C !B A)+(!D C B !A)+(!D C B A)), LSE_LINE_FILE_ID=3, LSE_LCOL=13, LSE_RCOL=44, LSE_LLINE=32, LSE_RLINE=32 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(11[2:53])
    defparam I1.init = 16'b0000000011111111;
    
endmodule
//
// Verilog Description of module inverter_U614
//

module inverter_U614 (\notGate[445]_keep , \notGate[446] ) /* synthesis syn_module_defined=1 */ ;
    input \notGate[445]_keep ;
    output \notGate[446] ;
    
    wire \notGate[445]_keep  /* synthesis alspreserve=1 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(25[15:22])
    
    LUT4 I1 (.A(\notGate[445]_keep ), .B(\notGate[445]_keep ), .C(\notGate[445]_keep ), 
         .D(\notGate[445]_keep ), .Z(\notGate[446] )) /* synthesis syn_instantiated=1, lut_function=((!D !C !B !A)+(!D !C !B A)+(!D !C B !A)+(!D !C B A)+(!D C !B !A)+(!D C !B A)+(!D C B !A)+(!D C B A)), LSE_LINE_FILE_ID=3, LSE_LCOL=13, LSE_RCOL=44, LSE_LLINE=32, LSE_RLINE=32 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(11[2:53])
    defparam I1.init = 16'b0000000011111111;
    
endmodule
//
// Verilog Description of module inverter_U615
//

module inverter_U615 (\notGate[444]_keep , \notGate[445] ) /* synthesis syn_module_defined=1 */ ;
    input \notGate[444]_keep ;
    output \notGate[445] ;
    
    wire \notGate[444]_keep  /* synthesis alspreserve=1 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(25[15:22])
    
    LUT4 I1 (.A(\notGate[444]_keep ), .B(\notGate[444]_keep ), .C(\notGate[444]_keep ), 
         .D(\notGate[444]_keep ), .Z(\notGate[445] )) /* synthesis syn_instantiated=1, lut_function=((!D !C !B !A)+(!D !C !B A)+(!D !C B !A)+(!D !C B A)+(!D C !B !A)+(!D C !B A)+(!D C B !A)+(!D C B A)), LSE_LINE_FILE_ID=3, LSE_LCOL=13, LSE_RCOL=44, LSE_LLINE=32, LSE_RLINE=32 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(11[2:53])
    defparam I1.init = 16'b0000000011111111;
    
endmodule
//
// Verilog Description of module inverter_U616
//

module inverter_U616 (\notGate[443]_keep , \notGate[444] ) /* synthesis syn_module_defined=1 */ ;
    input \notGate[443]_keep ;
    output \notGate[444] ;
    
    wire \notGate[443]_keep  /* synthesis alspreserve=1 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(25[15:22])
    
    LUT4 I1 (.A(\notGate[443]_keep ), .B(\notGate[443]_keep ), .C(\notGate[443]_keep ), 
         .D(\notGate[443]_keep ), .Z(\notGate[444] )) /* synthesis syn_instantiated=1, lut_function=((!D !C !B !A)+(!D !C !B A)+(!D !C B !A)+(!D !C B A)+(!D C !B !A)+(!D C !B A)+(!D C B !A)+(!D C B A)), LSE_LINE_FILE_ID=3, LSE_LCOL=13, LSE_RCOL=44, LSE_LLINE=32, LSE_RLINE=32 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(11[2:53])
    defparam I1.init = 16'b0000000011111111;
    
endmodule
//
// Verilog Description of module inverter_U617
//

module inverter_U617 (\notGate[442]_keep , \notGate[443] ) /* synthesis syn_module_defined=1 */ ;
    input \notGate[442]_keep ;
    output \notGate[443] ;
    
    wire \notGate[442]_keep  /* synthesis alspreserve=1 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(25[15:22])
    
    LUT4 I1 (.A(\notGate[442]_keep ), .B(\notGate[442]_keep ), .C(\notGate[442]_keep ), 
         .D(\notGate[442]_keep ), .Z(\notGate[443] )) /* synthesis syn_instantiated=1, lut_function=((!D !C !B !A)+(!D !C !B A)+(!D !C B !A)+(!D !C B A)+(!D C !B !A)+(!D C !B A)+(!D C B !A)+(!D C B A)), LSE_LINE_FILE_ID=3, LSE_LCOL=13, LSE_RCOL=44, LSE_LLINE=32, LSE_RLINE=32 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(11[2:53])
    defparam I1.init = 16'b0000000011111111;
    
endmodule
//
// Verilog Description of module inverter_U618
//

module inverter_U618 (\notGate[441]_keep , \notGate[442] ) /* synthesis syn_module_defined=1 */ ;
    input \notGate[441]_keep ;
    output \notGate[442] ;
    
    wire \notGate[441]_keep  /* synthesis alspreserve=1 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(25[15:22])
    
    LUT4 I1 (.A(\notGate[441]_keep ), .B(\notGate[441]_keep ), .C(\notGate[441]_keep ), 
         .D(\notGate[441]_keep ), .Z(\notGate[442] )) /* synthesis syn_instantiated=1, lut_function=((!D !C !B !A)+(!D !C !B A)+(!D !C B !A)+(!D !C B A)+(!D C !B !A)+(!D C !B A)+(!D C B !A)+(!D C B A)), LSE_LINE_FILE_ID=3, LSE_LCOL=13, LSE_RCOL=44, LSE_LLINE=32, LSE_RLINE=32 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(11[2:53])
    defparam I1.init = 16'b0000000011111111;
    
endmodule
//
// Verilog Description of module inverter_U619
//

module inverter_U619 (\notGate[440]_keep , \notGate[441] ) /* synthesis syn_module_defined=1 */ ;
    input \notGate[440]_keep ;
    output \notGate[441] ;
    
    wire \notGate[440]_keep  /* synthesis alspreserve=1 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(25[15:22])
    
    LUT4 I1 (.A(\notGate[440]_keep ), .B(\notGate[440]_keep ), .C(\notGate[440]_keep ), 
         .D(\notGate[440]_keep ), .Z(\notGate[441] )) /* synthesis syn_instantiated=1, lut_function=((!D !C !B !A)+(!D !C !B A)+(!D !C B !A)+(!D !C B A)+(!D C !B !A)+(!D C !B A)+(!D C B !A)+(!D C B A)), LSE_LINE_FILE_ID=3, LSE_LCOL=13, LSE_RCOL=44, LSE_LLINE=32, LSE_RLINE=32 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(11[2:53])
    defparam I1.init = 16'b0000000011111111;
    
endmodule
//
// Verilog Description of module inverter_U620
//

module inverter_U620 (\notGate[439]_keep , \notGate[440] ) /* synthesis syn_module_defined=1 */ ;
    input \notGate[439]_keep ;
    output \notGate[440] ;
    
    wire \notGate[439]_keep  /* synthesis alspreserve=1 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(25[15:22])
    
    LUT4 I1 (.A(\notGate[439]_keep ), .B(\notGate[439]_keep ), .C(\notGate[439]_keep ), 
         .D(\notGate[439]_keep ), .Z(\notGate[440] )) /* synthesis syn_instantiated=1, lut_function=((!D !C !B !A)+(!D !C !B A)+(!D !C B !A)+(!D !C B A)+(!D C !B !A)+(!D C !B A)+(!D C B !A)+(!D C B A)), LSE_LINE_FILE_ID=3, LSE_LCOL=13, LSE_RCOL=44, LSE_LLINE=32, LSE_RLINE=32 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(11[2:53])
    defparam I1.init = 16'b0000000011111111;
    
endmodule
//
// Verilog Description of module inverter_U621
//

module inverter_U621 (\notGate[42]_keep , \notGate[43] ) /* synthesis syn_module_defined=1 */ ;
    input \notGate[42]_keep ;
    output \notGate[43] ;
    
    wire \notGate[42]_keep  /* synthesis alspreserve=1 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(25[15:22])
    
    LUT4 I1 (.A(\notGate[42]_keep ), .B(\notGate[42]_keep ), .C(\notGate[42]_keep ), 
         .D(\notGate[42]_keep ), .Z(\notGate[43] )) /* synthesis syn_instantiated=1, lut_function=((!D !C !B !A)+(!D !C !B A)+(!D !C B !A)+(!D !C B A)+(!D C !B !A)+(!D C !B A)+(!D C B !A)+(!D C B A)), LSE_LINE_FILE_ID=3, LSE_LCOL=13, LSE_RCOL=44, LSE_LLINE=32, LSE_RLINE=32 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(11[2:53])
    defparam I1.init = 16'b0000000011111111;
    
endmodule
//
// Verilog Description of module inverter_U622
//

module inverter_U622 (\notGate[438]_keep , \notGate[439] ) /* synthesis syn_module_defined=1 */ ;
    input \notGate[438]_keep ;
    output \notGate[439] ;
    
    wire \notGate[438]_keep  /* synthesis alspreserve=1 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(25[15:22])
    
    LUT4 I1 (.A(\notGate[438]_keep ), .B(\notGate[438]_keep ), .C(\notGate[438]_keep ), 
         .D(\notGate[438]_keep ), .Z(\notGate[439] )) /* synthesis syn_instantiated=1, lut_function=((!D !C !B !A)+(!D !C !B A)+(!D !C B !A)+(!D !C B A)+(!D C !B !A)+(!D C !B A)+(!D C B !A)+(!D C B A)), LSE_LINE_FILE_ID=3, LSE_LCOL=13, LSE_RCOL=44, LSE_LLINE=32, LSE_RLINE=32 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(11[2:53])
    defparam I1.init = 16'b0000000011111111;
    
endmodule
//
// Verilog Description of module inverter_U623
//

module inverter_U623 (\notGate[437]_keep , \notGate[438] ) /* synthesis syn_module_defined=1 */ ;
    input \notGate[437]_keep ;
    output \notGate[438] ;
    
    wire \notGate[437]_keep  /* synthesis alspreserve=1 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(25[15:22])
    
    LUT4 I1 (.A(\notGate[437]_keep ), .B(\notGate[437]_keep ), .C(\notGate[437]_keep ), 
         .D(\notGate[437]_keep ), .Z(\notGate[438] )) /* synthesis syn_instantiated=1, lut_function=((!D !C !B !A)+(!D !C !B A)+(!D !C B !A)+(!D !C B A)+(!D C !B !A)+(!D C !B A)+(!D C B !A)+(!D C B A)), LSE_LINE_FILE_ID=3, LSE_LCOL=13, LSE_RCOL=44, LSE_LLINE=32, LSE_RLINE=32 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(11[2:53])
    defparam I1.init = 16'b0000000011111111;
    
endmodule
//
// Verilog Description of module inverter_U624
//

module inverter_U624 (\notGate[436]_keep , \notGate[437] ) /* synthesis syn_module_defined=1 */ ;
    input \notGate[436]_keep ;
    output \notGate[437] ;
    
    wire \notGate[436]_keep  /* synthesis alspreserve=1 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(25[15:22])
    
    LUT4 I1 (.A(\notGate[436]_keep ), .B(\notGate[436]_keep ), .C(\notGate[436]_keep ), 
         .D(\notGate[436]_keep ), .Z(\notGate[437] )) /* synthesis syn_instantiated=1, lut_function=((!D !C !B !A)+(!D !C !B A)+(!D !C B !A)+(!D !C B A)+(!D C !B !A)+(!D C !B A)+(!D C B !A)+(!D C B A)), LSE_LINE_FILE_ID=3, LSE_LCOL=13, LSE_RCOL=44, LSE_LLINE=32, LSE_RLINE=32 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(11[2:53])
    defparam I1.init = 16'b0000000011111111;
    
endmodule
//
// Verilog Description of module inverter_U625
//

module inverter_U625 (\notGate[435]_keep , \notGate[436] ) /* synthesis syn_module_defined=1 */ ;
    input \notGate[435]_keep ;
    output \notGate[436] ;
    
    wire \notGate[435]_keep  /* synthesis alspreserve=1 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(25[15:22])
    
    LUT4 I1 (.A(\notGate[435]_keep ), .B(\notGate[435]_keep ), .C(\notGate[435]_keep ), 
         .D(\notGate[435]_keep ), .Z(\notGate[436] )) /* synthesis syn_instantiated=1, lut_function=((!D !C !B !A)+(!D !C !B A)+(!D !C B !A)+(!D !C B A)+(!D C !B !A)+(!D C !B A)+(!D C B !A)+(!D C B A)), LSE_LINE_FILE_ID=3, LSE_LCOL=13, LSE_RCOL=44, LSE_LLINE=32, LSE_RLINE=32 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(11[2:53])
    defparam I1.init = 16'b0000000011111111;
    
endmodule
//
// Verilog Description of module inverter_U626
//

module inverter_U626 (\notGate[434]_keep , \notGate[435] ) /* synthesis syn_module_defined=1 */ ;
    input \notGate[434]_keep ;
    output \notGate[435] ;
    
    wire \notGate[434]_keep  /* synthesis alspreserve=1 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(25[15:22])
    
    LUT4 I1 (.A(\notGate[434]_keep ), .B(\notGate[434]_keep ), .C(\notGate[434]_keep ), 
         .D(\notGate[434]_keep ), .Z(\notGate[435] )) /* synthesis syn_instantiated=1, lut_function=((!D !C !B !A)+(!D !C !B A)+(!D !C B !A)+(!D !C B A)+(!D C !B !A)+(!D C !B A)+(!D C B !A)+(!D C B A)), LSE_LINE_FILE_ID=3, LSE_LCOL=13, LSE_RCOL=44, LSE_LLINE=32, LSE_RLINE=32 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(11[2:53])
    defparam I1.init = 16'b0000000011111111;
    
endmodule
//
// Verilog Description of module inverter_U627
//

module inverter_U627 (\notGate[433]_keep , \notGate[434] ) /* synthesis syn_module_defined=1 */ ;
    input \notGate[433]_keep ;
    output \notGate[434] ;
    
    wire \notGate[433]_keep  /* synthesis alspreserve=1 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(25[15:22])
    
    LUT4 I1 (.A(\notGate[433]_keep ), .B(\notGate[433]_keep ), .C(\notGate[433]_keep ), 
         .D(\notGate[433]_keep ), .Z(\notGate[434] )) /* synthesis syn_instantiated=1, lut_function=((!D !C !B !A)+(!D !C !B A)+(!D !C B !A)+(!D !C B A)+(!D C !B !A)+(!D C !B A)+(!D C B !A)+(!D C B A)), LSE_LINE_FILE_ID=3, LSE_LCOL=13, LSE_RCOL=44, LSE_LLINE=32, LSE_RLINE=32 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(11[2:53])
    defparam I1.init = 16'b0000000011111111;
    
endmodule
//
// Verilog Description of module inverter_U628
//

module inverter_U628 (\notGate[432]_keep , \notGate[433] ) /* synthesis syn_module_defined=1 */ ;
    input \notGate[432]_keep ;
    output \notGate[433] ;
    
    wire \notGate[432]_keep  /* synthesis alspreserve=1 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(25[15:22])
    
    LUT4 I1 (.A(\notGate[432]_keep ), .B(\notGate[432]_keep ), .C(\notGate[432]_keep ), 
         .D(\notGate[432]_keep ), .Z(\notGate[433] )) /* synthesis syn_instantiated=1, lut_function=((!D !C !B !A)+(!D !C !B A)+(!D !C B !A)+(!D !C B A)+(!D C !B !A)+(!D C !B A)+(!D C B !A)+(!D C B A)), LSE_LINE_FILE_ID=3, LSE_LCOL=13, LSE_RCOL=44, LSE_LLINE=32, LSE_RLINE=32 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(11[2:53])
    defparam I1.init = 16'b0000000011111111;
    
endmodule
//
// Verilog Description of module inverter_U629
//

module inverter_U629 (\notGate[431]_keep , \notGate[432] ) /* synthesis syn_module_defined=1 */ ;
    input \notGate[431]_keep ;
    output \notGate[432] ;
    
    wire \notGate[431]_keep  /* synthesis alspreserve=1 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(25[15:22])
    
    LUT4 I1 (.A(\notGate[431]_keep ), .B(\notGate[431]_keep ), .C(\notGate[431]_keep ), 
         .D(\notGate[431]_keep ), .Z(\notGate[432] )) /* synthesis syn_instantiated=1, lut_function=((!D !C !B !A)+(!D !C !B A)+(!D !C B !A)+(!D !C B A)+(!D C !B !A)+(!D C !B A)+(!D C B !A)+(!D C B A)), LSE_LINE_FILE_ID=3, LSE_LCOL=13, LSE_RCOL=44, LSE_LLINE=32, LSE_RLINE=32 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(11[2:53])
    defparam I1.init = 16'b0000000011111111;
    
endmodule
//
// Verilog Description of module inverter_U630
//

module inverter_U630 (\notGate[430]_keep , \notGate[431] ) /* synthesis syn_module_defined=1 */ ;
    input \notGate[430]_keep ;
    output \notGate[431] ;
    
    wire \notGate[430]_keep  /* synthesis alspreserve=1 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(25[15:22])
    
    LUT4 I1 (.A(\notGate[430]_keep ), .B(\notGate[430]_keep ), .C(\notGate[430]_keep ), 
         .D(\notGate[430]_keep ), .Z(\notGate[431] )) /* synthesis syn_instantiated=1, lut_function=((!D !C !B !A)+(!D !C !B A)+(!D !C B !A)+(!D !C B A)+(!D C !B !A)+(!D C !B A)+(!D C B !A)+(!D C B A)), LSE_LINE_FILE_ID=3, LSE_LCOL=13, LSE_RCOL=44, LSE_LLINE=32, LSE_RLINE=32 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(11[2:53])
    defparam I1.init = 16'b0000000011111111;
    
endmodule
//
// Verilog Description of module inverter_U631
//

module inverter_U631 (\notGate[429]_keep , \notGate[430] ) /* synthesis syn_module_defined=1 */ ;
    input \notGate[429]_keep ;
    output \notGate[430] ;
    
    wire \notGate[429]_keep  /* synthesis alspreserve=1 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(25[15:22])
    
    LUT4 I1 (.A(\notGate[429]_keep ), .B(\notGate[429]_keep ), .C(\notGate[429]_keep ), 
         .D(\notGate[429]_keep ), .Z(\notGate[430] )) /* synthesis syn_instantiated=1, lut_function=((!D !C !B !A)+(!D !C !B A)+(!D !C B !A)+(!D !C B A)+(!D C !B !A)+(!D C !B A)+(!D C B !A)+(!D C B A)), LSE_LINE_FILE_ID=3, LSE_LCOL=13, LSE_RCOL=44, LSE_LLINE=32, LSE_RLINE=32 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(11[2:53])
    defparam I1.init = 16'b0000000011111111;
    
endmodule
//
// Verilog Description of module inverter_U632
//

module inverter_U632 (\notGate[41]_keep , \notGate[42] ) /* synthesis syn_module_defined=1 */ ;
    input \notGate[41]_keep ;
    output \notGate[42] ;
    
    wire \notGate[41]_keep  /* synthesis alspreserve=1 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(25[15:22])
    
    LUT4 I1 (.A(\notGate[41]_keep ), .B(\notGate[41]_keep ), .C(\notGate[41]_keep ), 
         .D(\notGate[41]_keep ), .Z(\notGate[42] )) /* synthesis syn_instantiated=1, lut_function=((!D !C !B !A)+(!D !C !B A)+(!D !C B !A)+(!D !C B A)+(!D C !B !A)+(!D C !B A)+(!D C B !A)+(!D C B A)), LSE_LINE_FILE_ID=3, LSE_LCOL=13, LSE_RCOL=44, LSE_LLINE=32, LSE_RLINE=32 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(11[2:53])
    defparam I1.init = 16'b0000000011111111;
    
endmodule
//
// Verilog Description of module inverter_U633
//

module inverter_U633 (\notGate[428]_keep , \notGate[429] ) /* synthesis syn_module_defined=1 */ ;
    input \notGate[428]_keep ;
    output \notGate[429] ;
    
    wire \notGate[428]_keep  /* synthesis alspreserve=1 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(25[15:22])
    
    LUT4 I1 (.A(\notGate[428]_keep ), .B(\notGate[428]_keep ), .C(\notGate[428]_keep ), 
         .D(\notGate[428]_keep ), .Z(\notGate[429] )) /* synthesis syn_instantiated=1, lut_function=((!D !C !B !A)+(!D !C !B A)+(!D !C B !A)+(!D !C B A)+(!D C !B !A)+(!D C !B A)+(!D C B !A)+(!D C B A)), LSE_LINE_FILE_ID=3, LSE_LCOL=13, LSE_RCOL=44, LSE_LLINE=32, LSE_RLINE=32 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(11[2:53])
    defparam I1.init = 16'b0000000011111111;
    
endmodule
//
// Verilog Description of module inverter_U634
//

module inverter_U634 (\notGate[427]_keep , \notGate[428] ) /* synthesis syn_module_defined=1 */ ;
    input \notGate[427]_keep ;
    output \notGate[428] ;
    
    wire \notGate[427]_keep  /* synthesis alspreserve=1 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(25[15:22])
    
    LUT4 I1 (.A(\notGate[427]_keep ), .B(\notGate[427]_keep ), .C(\notGate[427]_keep ), 
         .D(\notGate[427]_keep ), .Z(\notGate[428] )) /* synthesis syn_instantiated=1, lut_function=((!D !C !B !A)+(!D !C !B A)+(!D !C B !A)+(!D !C B A)+(!D C !B !A)+(!D C !B A)+(!D C B !A)+(!D C B A)), LSE_LINE_FILE_ID=3, LSE_LCOL=13, LSE_RCOL=44, LSE_LLINE=32, LSE_RLINE=32 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(11[2:53])
    defparam I1.init = 16'b0000000011111111;
    
endmodule
//
// Verilog Description of module inverter_U635
//

module inverter_U635 (\notGate[426]_keep , \notGate[427] ) /* synthesis syn_module_defined=1 */ ;
    input \notGate[426]_keep ;
    output \notGate[427] ;
    
    wire \notGate[426]_keep  /* synthesis alspreserve=1 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(25[15:22])
    
    LUT4 I1 (.A(\notGate[426]_keep ), .B(\notGate[426]_keep ), .C(\notGate[426]_keep ), 
         .D(\notGate[426]_keep ), .Z(\notGate[427] )) /* synthesis syn_instantiated=1, lut_function=((!D !C !B !A)+(!D !C !B A)+(!D !C B !A)+(!D !C B A)+(!D C !B !A)+(!D C !B A)+(!D C B !A)+(!D C B A)), LSE_LINE_FILE_ID=3, LSE_LCOL=13, LSE_RCOL=44, LSE_LLINE=32, LSE_RLINE=32 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(11[2:53])
    defparam I1.init = 16'b0000000011111111;
    
endmodule
//
// Verilog Description of module inverter_U636
//

module inverter_U636 (\notGate[425]_keep , \notGate[426] ) /* synthesis syn_module_defined=1 */ ;
    input \notGate[425]_keep ;
    output \notGate[426] ;
    
    wire \notGate[425]_keep  /* synthesis alspreserve=1 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(25[15:22])
    
    LUT4 I1 (.A(\notGate[425]_keep ), .B(\notGate[425]_keep ), .C(\notGate[425]_keep ), 
         .D(\notGate[425]_keep ), .Z(\notGate[426] )) /* synthesis syn_instantiated=1, lut_function=((!D !C !B !A)+(!D !C !B A)+(!D !C B !A)+(!D !C B A)+(!D C !B !A)+(!D C !B A)+(!D C B !A)+(!D C B A)), LSE_LINE_FILE_ID=3, LSE_LCOL=13, LSE_RCOL=44, LSE_LLINE=32, LSE_RLINE=32 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(11[2:53])
    defparam I1.init = 16'b0000000011111111;
    
endmodule
//
// Verilog Description of module inverter_U637
//

module inverter_U637 (\notGate[424]_keep , \notGate[425] ) /* synthesis syn_module_defined=1 */ ;
    input \notGate[424]_keep ;
    output \notGate[425] ;
    
    wire \notGate[424]_keep  /* synthesis alspreserve=1 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(25[15:22])
    
    LUT4 I1 (.A(\notGate[424]_keep ), .B(\notGate[424]_keep ), .C(\notGate[424]_keep ), 
         .D(\notGate[424]_keep ), .Z(\notGate[425] )) /* synthesis syn_instantiated=1, lut_function=((!D !C !B !A)+(!D !C !B A)+(!D !C B !A)+(!D !C B A)+(!D C !B !A)+(!D C !B A)+(!D C B !A)+(!D C B A)), LSE_LINE_FILE_ID=3, LSE_LCOL=13, LSE_RCOL=44, LSE_LLINE=32, LSE_RLINE=32 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(11[2:53])
    defparam I1.init = 16'b0000000011111111;
    
endmodule
//
// Verilog Description of module inverter_U638
//

module inverter_U638 (\notGate[423]_keep , \notGate[424] ) /* synthesis syn_module_defined=1 */ ;
    input \notGate[423]_keep ;
    output \notGate[424] ;
    
    wire \notGate[423]_keep  /* synthesis alspreserve=1 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(25[15:22])
    
    LUT4 I1 (.A(\notGate[423]_keep ), .B(\notGate[423]_keep ), .C(\notGate[423]_keep ), 
         .D(\notGate[423]_keep ), .Z(\notGate[424] )) /* synthesis syn_instantiated=1, lut_function=((!D !C !B !A)+(!D !C !B A)+(!D !C B !A)+(!D !C B A)+(!D C !B !A)+(!D C !B A)+(!D C B !A)+(!D C B A)), LSE_LINE_FILE_ID=3, LSE_LCOL=13, LSE_RCOL=44, LSE_LLINE=32, LSE_RLINE=32 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(11[2:53])
    defparam I1.init = 16'b0000000011111111;
    
endmodule
//
// Verilog Description of module inverter_U639
//

module inverter_U639 (\notGate[422]_keep , \notGate[423] ) /* synthesis syn_module_defined=1 */ ;
    input \notGate[422]_keep ;
    output \notGate[423] ;
    
    wire \notGate[422]_keep  /* synthesis alspreserve=1 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(25[15:22])
    
    LUT4 I1 (.A(\notGate[422]_keep ), .B(\notGate[422]_keep ), .C(\notGate[422]_keep ), 
         .D(\notGate[422]_keep ), .Z(\notGate[423] )) /* synthesis syn_instantiated=1, lut_function=((!D !C !B !A)+(!D !C !B A)+(!D !C B !A)+(!D !C B A)+(!D C !B !A)+(!D C !B A)+(!D C B !A)+(!D C B A)), LSE_LINE_FILE_ID=3, LSE_LCOL=13, LSE_RCOL=44, LSE_LLINE=32, LSE_RLINE=32 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(11[2:53])
    defparam I1.init = 16'b0000000011111111;
    
endmodule
//
// Verilog Description of module inverter_U640
//

module inverter_U640 (\notGate[421]_keep , \notGate[422] ) /* synthesis syn_module_defined=1 */ ;
    input \notGate[421]_keep ;
    output \notGate[422] ;
    
    wire \notGate[421]_keep  /* synthesis alspreserve=1 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(25[15:22])
    
    LUT4 I1 (.A(\notGate[421]_keep ), .B(\notGate[421]_keep ), .C(\notGate[421]_keep ), 
         .D(\notGate[421]_keep ), .Z(\notGate[422] )) /* synthesis syn_instantiated=1, lut_function=((!D !C !B !A)+(!D !C !B A)+(!D !C B !A)+(!D !C B A)+(!D C !B !A)+(!D C !B A)+(!D C B !A)+(!D C B A)), LSE_LINE_FILE_ID=3, LSE_LCOL=13, LSE_RCOL=44, LSE_LLINE=32, LSE_RLINE=32 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(11[2:53])
    defparam I1.init = 16'b0000000011111111;
    
endmodule
//
// Verilog Description of module inverter_U641
//

module inverter_U641 (\notGate[420]_keep , \notGate[421] ) /* synthesis syn_module_defined=1 */ ;
    input \notGate[420]_keep ;
    output \notGate[421] ;
    
    wire \notGate[420]_keep  /* synthesis alspreserve=1 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(25[15:22])
    
    LUT4 I1 (.A(\notGate[420]_keep ), .B(\notGate[420]_keep ), .C(\notGate[420]_keep ), 
         .D(\notGate[420]_keep ), .Z(\notGate[421] )) /* synthesis syn_instantiated=1, lut_function=((!D !C !B !A)+(!D !C !B A)+(!D !C B !A)+(!D !C B A)+(!D C !B !A)+(!D C !B A)+(!D C B !A)+(!D C B A)), LSE_LINE_FILE_ID=3, LSE_LCOL=13, LSE_RCOL=44, LSE_LLINE=32, LSE_RLINE=32 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(11[2:53])
    defparam I1.init = 16'b0000000011111111;
    
endmodule
//
// Verilog Description of module inverter_U642
//

module inverter_U642 (\notGate[419]_keep , \notGate[420] ) /* synthesis syn_module_defined=1 */ ;
    input \notGate[419]_keep ;
    output \notGate[420] ;
    
    wire \notGate[419]_keep  /* synthesis alspreserve=1 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(25[15:22])
    
    LUT4 I1 (.A(\notGate[419]_keep ), .B(\notGate[419]_keep ), .C(\notGate[419]_keep ), 
         .D(\notGate[419]_keep ), .Z(\notGate[420] )) /* synthesis syn_instantiated=1, lut_function=((!D !C !B !A)+(!D !C !B A)+(!D !C B !A)+(!D !C B A)+(!D C !B !A)+(!D C !B A)+(!D C B !A)+(!D C B A)), LSE_LINE_FILE_ID=3, LSE_LCOL=13, LSE_RCOL=44, LSE_LLINE=32, LSE_RLINE=32 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(11[2:53])
    defparam I1.init = 16'b0000000011111111;
    
endmodule
//
// Verilog Description of module inverter_U643
//

module inverter_U643 (\notGate[40]_keep , \notGate[41] ) /* synthesis syn_module_defined=1 */ ;
    input \notGate[40]_keep ;
    output \notGate[41] ;
    
    wire \notGate[40]_keep  /* synthesis alspreserve=1 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(25[15:22])
    
    LUT4 I1 (.A(\notGate[40]_keep ), .B(\notGate[40]_keep ), .C(\notGate[40]_keep ), 
         .D(\notGate[40]_keep ), .Z(\notGate[41] )) /* synthesis syn_instantiated=1, lut_function=((!D !C !B !A)+(!D !C !B A)+(!D !C B !A)+(!D !C B A)+(!D C !B !A)+(!D C !B A)+(!D C B !A)+(!D C B A)), LSE_LINE_FILE_ID=3, LSE_LCOL=13, LSE_RCOL=44, LSE_LLINE=32, LSE_RLINE=32 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(11[2:53])
    defparam I1.init = 16'b0000000011111111;
    
endmodule
//
// Verilog Description of module inverter_U644
//

module inverter_U644 (\notGate[418]_keep , \notGate[419] ) /* synthesis syn_module_defined=1 */ ;
    input \notGate[418]_keep ;
    output \notGate[419] ;
    
    wire \notGate[418]_keep  /* synthesis alspreserve=1 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(25[15:22])
    
    LUT4 I1 (.A(\notGate[418]_keep ), .B(\notGate[418]_keep ), .C(\notGate[418]_keep ), 
         .D(\notGate[418]_keep ), .Z(\notGate[419] )) /* synthesis syn_instantiated=1, lut_function=((!D !C !B !A)+(!D !C !B A)+(!D !C B !A)+(!D !C B A)+(!D C !B !A)+(!D C !B A)+(!D C B !A)+(!D C B A)), LSE_LINE_FILE_ID=3, LSE_LCOL=13, LSE_RCOL=44, LSE_LLINE=32, LSE_RLINE=32 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(11[2:53])
    defparam I1.init = 16'b0000000011111111;
    
endmodule
//
// Verilog Description of module inverter_U645
//

module inverter_U645 (\notGate[417]_keep , \notGate[418] ) /* synthesis syn_module_defined=1 */ ;
    input \notGate[417]_keep ;
    output \notGate[418] ;
    
    wire \notGate[417]_keep  /* synthesis alspreserve=1 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(25[15:22])
    
    LUT4 I1 (.A(\notGate[417]_keep ), .B(\notGate[417]_keep ), .C(\notGate[417]_keep ), 
         .D(\notGate[417]_keep ), .Z(\notGate[418] )) /* synthesis syn_instantiated=1, lut_function=((!D !C !B !A)+(!D !C !B A)+(!D !C B !A)+(!D !C B A)+(!D C !B !A)+(!D C !B A)+(!D C B !A)+(!D C B A)), LSE_LINE_FILE_ID=3, LSE_LCOL=13, LSE_RCOL=44, LSE_LLINE=32, LSE_RLINE=32 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(11[2:53])
    defparam I1.init = 16'b0000000011111111;
    
endmodule
//
// Verilog Description of module inverter_U646
//

module inverter_U646 (\notGate[416]_keep , \notGate[417] ) /* synthesis syn_module_defined=1 */ ;
    input \notGate[416]_keep ;
    output \notGate[417] ;
    
    wire \notGate[416]_keep  /* synthesis alspreserve=1 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(25[15:22])
    
    LUT4 I1 (.A(\notGate[416]_keep ), .B(\notGate[416]_keep ), .C(\notGate[416]_keep ), 
         .D(\notGate[416]_keep ), .Z(\notGate[417] )) /* synthesis syn_instantiated=1, lut_function=((!D !C !B !A)+(!D !C !B A)+(!D !C B !A)+(!D !C B A)+(!D C !B !A)+(!D C !B A)+(!D C B !A)+(!D C B A)), LSE_LINE_FILE_ID=3, LSE_LCOL=13, LSE_RCOL=44, LSE_LLINE=32, LSE_RLINE=32 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(11[2:53])
    defparam I1.init = 16'b0000000011111111;
    
endmodule
//
// Verilog Description of module inverter_U647
//

module inverter_U647 (\notGate[415]_keep , \notGate[416] ) /* synthesis syn_module_defined=1 */ ;
    input \notGate[415]_keep ;
    output \notGate[416] ;
    
    wire \notGate[415]_keep  /* synthesis alspreserve=1 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(25[15:22])
    
    LUT4 I1 (.A(\notGate[415]_keep ), .B(\notGate[415]_keep ), .C(\notGate[415]_keep ), 
         .D(\notGate[415]_keep ), .Z(\notGate[416] )) /* synthesis syn_instantiated=1, lut_function=((!D !C !B !A)+(!D !C !B A)+(!D !C B !A)+(!D !C B A)+(!D C !B !A)+(!D C !B A)+(!D C B !A)+(!D C B A)), LSE_LINE_FILE_ID=3, LSE_LCOL=13, LSE_RCOL=44, LSE_LLINE=32, LSE_RLINE=32 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(11[2:53])
    defparam I1.init = 16'b0000000011111111;
    
endmodule
//
// Verilog Description of module inverter_U648
//

module inverter_U648 (\notGate[414]_keep , \notGate[415] ) /* synthesis syn_module_defined=1 */ ;
    input \notGate[414]_keep ;
    output \notGate[415] ;
    
    wire \notGate[414]_keep  /* synthesis alspreserve=1 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(25[15:22])
    
    LUT4 I1 (.A(\notGate[414]_keep ), .B(\notGate[414]_keep ), .C(\notGate[414]_keep ), 
         .D(\notGate[414]_keep ), .Z(\notGate[415] )) /* synthesis syn_instantiated=1, lut_function=((!D !C !B !A)+(!D !C !B A)+(!D !C B !A)+(!D !C B A)+(!D C !B !A)+(!D C !B A)+(!D C B !A)+(!D C B A)), LSE_LINE_FILE_ID=3, LSE_LCOL=13, LSE_RCOL=44, LSE_LLINE=32, LSE_RLINE=32 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(11[2:53])
    defparam I1.init = 16'b0000000011111111;
    
endmodule
//
// Verilog Description of module inverter_U649
//

module inverter_U649 (\notGate[413]_keep , \notGate[414] ) /* synthesis syn_module_defined=1 */ ;
    input \notGate[413]_keep ;
    output \notGate[414] ;
    
    wire \notGate[413]_keep  /* synthesis alspreserve=1 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(25[15:22])
    
    LUT4 I1 (.A(\notGate[413]_keep ), .B(\notGate[413]_keep ), .C(\notGate[413]_keep ), 
         .D(\notGate[413]_keep ), .Z(\notGate[414] )) /* synthesis syn_instantiated=1, lut_function=((!D !C !B !A)+(!D !C !B A)+(!D !C B !A)+(!D !C B A)+(!D C !B !A)+(!D C !B A)+(!D C B !A)+(!D C B A)), LSE_LINE_FILE_ID=3, LSE_LCOL=13, LSE_RCOL=44, LSE_LLINE=32, LSE_RLINE=32 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(11[2:53])
    defparam I1.init = 16'b0000000011111111;
    
endmodule
//
// Verilog Description of module inverter_U650
//

module inverter_U650 (\notGate[412]_keep , \notGate[413] ) /* synthesis syn_module_defined=1 */ ;
    input \notGate[412]_keep ;
    output \notGate[413] ;
    
    wire \notGate[412]_keep  /* synthesis alspreserve=1 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(25[15:22])
    
    LUT4 I1 (.A(\notGate[412]_keep ), .B(\notGate[412]_keep ), .C(\notGate[412]_keep ), 
         .D(\notGate[412]_keep ), .Z(\notGate[413] )) /* synthesis syn_instantiated=1, lut_function=((!D !C !B !A)+(!D !C !B A)+(!D !C B !A)+(!D !C B A)+(!D C !B !A)+(!D C !B A)+(!D C B !A)+(!D C B A)), LSE_LINE_FILE_ID=3, LSE_LCOL=13, LSE_RCOL=44, LSE_LLINE=32, LSE_RLINE=32 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(11[2:53])
    defparam I1.init = 16'b0000000011111111;
    
endmodule
//
// Verilog Description of module inverter_U651
//

module inverter_U651 (\notGate[411]_keep , \notGate[412] ) /* synthesis syn_module_defined=1 */ ;
    input \notGate[411]_keep ;
    output \notGate[412] ;
    
    wire \notGate[411]_keep  /* synthesis alspreserve=1 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(25[15:22])
    
    LUT4 I1 (.A(\notGate[411]_keep ), .B(\notGate[411]_keep ), .C(\notGate[411]_keep ), 
         .D(\notGate[411]_keep ), .Z(\notGate[412] )) /* synthesis syn_instantiated=1, lut_function=((!D !C !B !A)+(!D !C !B A)+(!D !C B !A)+(!D !C B A)+(!D C !B !A)+(!D C !B A)+(!D C B !A)+(!D C B A)), LSE_LINE_FILE_ID=3, LSE_LCOL=13, LSE_RCOL=44, LSE_LLINE=32, LSE_RLINE=32 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(11[2:53])
    defparam I1.init = 16'b0000000011111111;
    
endmodule
//
// Verilog Description of module inverter_U652
//

module inverter_U652 (\notGate[410]_keep , \notGate[411] ) /* synthesis syn_module_defined=1 */ ;
    input \notGate[410]_keep ;
    output \notGate[411] ;
    
    wire \notGate[410]_keep  /* synthesis alspreserve=1 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(25[15:22])
    
    LUT4 I1 (.A(\notGate[410]_keep ), .B(\notGate[410]_keep ), .C(\notGate[410]_keep ), 
         .D(\notGate[410]_keep ), .Z(\notGate[411] )) /* synthesis syn_instantiated=1, lut_function=((!D !C !B !A)+(!D !C !B A)+(!D !C B !A)+(!D !C B A)+(!D C !B !A)+(!D C !B A)+(!D C B !A)+(!D C B A)), LSE_LINE_FILE_ID=3, LSE_LCOL=13, LSE_RCOL=44, LSE_LLINE=32, LSE_RLINE=32 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(11[2:53])
    defparam I1.init = 16'b0000000011111111;
    
endmodule
//
// Verilog Description of module inverter_U653
//

module inverter_U653 (\notGate[409]_keep , \notGate[410] ) /* synthesis syn_module_defined=1 */ ;
    input \notGate[409]_keep ;
    output \notGate[410] ;
    
    wire \notGate[409]_keep  /* synthesis alspreserve=1 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(25[15:22])
    
    LUT4 I1 (.A(\notGate[409]_keep ), .B(\notGate[409]_keep ), .C(\notGate[409]_keep ), 
         .D(\notGate[409]_keep ), .Z(\notGate[410] )) /* synthesis syn_instantiated=1, lut_function=((!D !C !B !A)+(!D !C !B A)+(!D !C B !A)+(!D !C B A)+(!D C !B !A)+(!D C !B A)+(!D C B !A)+(!D C B A)), LSE_LINE_FILE_ID=3, LSE_LCOL=13, LSE_RCOL=44, LSE_LLINE=32, LSE_RLINE=32 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(11[2:53])
    defparam I1.init = 16'b0000000011111111;
    
endmodule
//
// Verilog Description of module inverter_U654
//

module inverter_U654 (\notGate[39]_keep , \notGate[40] ) /* synthesis syn_module_defined=1 */ ;
    input \notGate[39]_keep ;
    output \notGate[40] ;
    
    wire \notGate[39]_keep  /* synthesis alspreserve=1 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(25[15:22])
    
    LUT4 I1 (.A(\notGate[39]_keep ), .B(\notGate[39]_keep ), .C(\notGate[39]_keep ), 
         .D(\notGate[39]_keep ), .Z(\notGate[40] )) /* synthesis syn_instantiated=1, lut_function=((!D !C !B !A)+(!D !C !B A)+(!D !C B !A)+(!D !C B A)+(!D C !B !A)+(!D C !B A)+(!D C B !A)+(!D C B A)), LSE_LINE_FILE_ID=3, LSE_LCOL=13, LSE_RCOL=44, LSE_LLINE=32, LSE_RLINE=32 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(11[2:53])
    defparam I1.init = 16'b0000000011111111;
    
endmodule
//
// Verilog Description of module inverter_U655
//

module inverter_U655 (\notGate[408]_keep , \notGate[409] ) /* synthesis syn_module_defined=1 */ ;
    input \notGate[408]_keep ;
    output \notGate[409] ;
    
    wire \notGate[408]_keep  /* synthesis alspreserve=1 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(25[15:22])
    
    LUT4 I1 (.A(\notGate[408]_keep ), .B(\notGate[408]_keep ), .C(\notGate[408]_keep ), 
         .D(\notGate[408]_keep ), .Z(\notGate[409] )) /* synthesis syn_instantiated=1, lut_function=((!D !C !B !A)+(!D !C !B A)+(!D !C B !A)+(!D !C B A)+(!D C !B !A)+(!D C !B A)+(!D C B !A)+(!D C B A)), LSE_LINE_FILE_ID=3, LSE_LCOL=13, LSE_RCOL=44, LSE_LLINE=32, LSE_RLINE=32 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(11[2:53])
    defparam I1.init = 16'b0000000011111111;
    
endmodule
//
// Verilog Description of module inverter_U656
//

module inverter_U656 (\notGate[407]_keep , \notGate[408] ) /* synthesis syn_module_defined=1 */ ;
    input \notGate[407]_keep ;
    output \notGate[408] ;
    
    wire \notGate[407]_keep  /* synthesis alspreserve=1 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(25[15:22])
    
    LUT4 I1 (.A(\notGate[407]_keep ), .B(\notGate[407]_keep ), .C(\notGate[407]_keep ), 
         .D(\notGate[407]_keep ), .Z(\notGate[408] )) /* synthesis syn_instantiated=1, lut_function=((!D !C !B !A)+(!D !C !B A)+(!D !C B !A)+(!D !C B A)+(!D C !B !A)+(!D C !B A)+(!D C B !A)+(!D C B A)), LSE_LINE_FILE_ID=3, LSE_LCOL=13, LSE_RCOL=44, LSE_LLINE=32, LSE_RLINE=32 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(11[2:53])
    defparam I1.init = 16'b0000000011111111;
    
endmodule
//
// Verilog Description of module inverter_U657
//

module inverter_U657 (\notGate[406]_keep , \notGate[407] ) /* synthesis syn_module_defined=1 */ ;
    input \notGate[406]_keep ;
    output \notGate[407] ;
    
    wire \notGate[406]_keep  /* synthesis alspreserve=1 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(25[15:22])
    
    LUT4 I1 (.A(\notGate[406]_keep ), .B(\notGate[406]_keep ), .C(\notGate[406]_keep ), 
         .D(\notGate[406]_keep ), .Z(\notGate[407] )) /* synthesis syn_instantiated=1, lut_function=((!D !C !B !A)+(!D !C !B A)+(!D !C B !A)+(!D !C B A)+(!D C !B !A)+(!D C !B A)+(!D C B !A)+(!D C B A)), LSE_LINE_FILE_ID=3, LSE_LCOL=13, LSE_RCOL=44, LSE_LLINE=32, LSE_RLINE=32 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(11[2:53])
    defparam I1.init = 16'b0000000011111111;
    
endmodule
//
// Verilog Description of module inverter_U658
//

module inverter_U658 (\notGate[405]_keep , \notGate[406] ) /* synthesis syn_module_defined=1 */ ;
    input \notGate[405]_keep ;
    output \notGate[406] ;
    
    wire \notGate[405]_keep  /* synthesis alspreserve=1 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(25[15:22])
    
    LUT4 I1 (.A(\notGate[405]_keep ), .B(\notGate[405]_keep ), .C(\notGate[405]_keep ), 
         .D(\notGate[405]_keep ), .Z(\notGate[406] )) /* synthesis syn_instantiated=1, lut_function=((!D !C !B !A)+(!D !C !B A)+(!D !C B !A)+(!D !C B A)+(!D C !B !A)+(!D C !B A)+(!D C B !A)+(!D C B A)), LSE_LINE_FILE_ID=3, LSE_LCOL=13, LSE_RCOL=44, LSE_LLINE=32, LSE_RLINE=32 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(11[2:53])
    defparam I1.init = 16'b0000000011111111;
    
endmodule
//
// Verilog Description of module inverter_U659
//

module inverter_U659 (\notGate[404]_keep , \notGate[405] ) /* synthesis syn_module_defined=1 */ ;
    input \notGate[404]_keep ;
    output \notGate[405] ;
    
    wire \notGate[404]_keep  /* synthesis alspreserve=1 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(25[15:22])
    
    LUT4 I1 (.A(\notGate[404]_keep ), .B(\notGate[404]_keep ), .C(\notGate[404]_keep ), 
         .D(\notGate[404]_keep ), .Z(\notGate[405] )) /* synthesis syn_instantiated=1, lut_function=((!D !C !B !A)+(!D !C !B A)+(!D !C B !A)+(!D !C B A)+(!D C !B !A)+(!D C !B A)+(!D C B !A)+(!D C B A)), LSE_LINE_FILE_ID=3, LSE_LCOL=13, LSE_RCOL=44, LSE_LLINE=32, LSE_RLINE=32 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(11[2:53])
    defparam I1.init = 16'b0000000011111111;
    
endmodule
//
// Verilog Description of module inverter_U660
//

module inverter_U660 (\notGate[403]_keep , \notGate[404] ) /* synthesis syn_module_defined=1 */ ;
    input \notGate[403]_keep ;
    output \notGate[404] ;
    
    wire \notGate[403]_keep  /* synthesis alspreserve=1 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(25[15:22])
    
    LUT4 I1 (.A(\notGate[403]_keep ), .B(\notGate[403]_keep ), .C(\notGate[403]_keep ), 
         .D(\notGate[403]_keep ), .Z(\notGate[404] )) /* synthesis syn_instantiated=1, lut_function=((!D !C !B !A)+(!D !C !B A)+(!D !C B !A)+(!D !C B A)+(!D C !B !A)+(!D C !B A)+(!D C B !A)+(!D C B A)), LSE_LINE_FILE_ID=3, LSE_LCOL=13, LSE_RCOL=44, LSE_LLINE=32, LSE_RLINE=32 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(11[2:53])
    defparam I1.init = 16'b0000000011111111;
    
endmodule
//
// Verilog Description of module inverter_U661
//

module inverter_U661 (\notGate[402]_keep , \notGate[403] ) /* synthesis syn_module_defined=1 */ ;
    input \notGate[402]_keep ;
    output \notGate[403] ;
    
    wire \notGate[402]_keep  /* synthesis alspreserve=1 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(25[15:22])
    
    LUT4 I1 (.A(\notGate[402]_keep ), .B(\notGate[402]_keep ), .C(\notGate[402]_keep ), 
         .D(\notGate[402]_keep ), .Z(\notGate[403] )) /* synthesis syn_instantiated=1, lut_function=((!D !C !B !A)+(!D !C !B A)+(!D !C B !A)+(!D !C B A)+(!D C !B !A)+(!D C !B A)+(!D C B !A)+(!D C B A)), LSE_LINE_FILE_ID=3, LSE_LCOL=13, LSE_RCOL=44, LSE_LLINE=32, LSE_RLINE=32 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(11[2:53])
    defparam I1.init = 16'b0000000011111111;
    
endmodule
//
// Verilog Description of module inverter_U662
//

module inverter_U662 (\notGate[401]_keep , \notGate[402] ) /* synthesis syn_module_defined=1 */ ;
    input \notGate[401]_keep ;
    output \notGate[402] ;
    
    wire \notGate[401]_keep  /* synthesis alspreserve=1 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(25[15:22])
    
    LUT4 I1 (.A(\notGate[401]_keep ), .B(\notGate[401]_keep ), .C(\notGate[401]_keep ), 
         .D(\notGate[401]_keep ), .Z(\notGate[402] )) /* synthesis syn_instantiated=1, lut_function=((!D !C !B !A)+(!D !C !B A)+(!D !C B !A)+(!D !C B A)+(!D C !B !A)+(!D C !B A)+(!D C B !A)+(!D C B A)), LSE_LINE_FILE_ID=3, LSE_LCOL=13, LSE_RCOL=44, LSE_LLINE=32, LSE_RLINE=32 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(11[2:53])
    defparam I1.init = 16'b0000000011111111;
    
endmodule
//
// Verilog Description of module inverter_U663
//

module inverter_U663 (\notGate[400]_keep , \notGate[401] ) /* synthesis syn_module_defined=1 */ ;
    input \notGate[400]_keep ;
    output \notGate[401] ;
    
    wire \notGate[400]_keep  /* synthesis alspreserve=1 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(25[15:22])
    
    LUT4 I1 (.A(\notGate[400]_keep ), .B(\notGate[400]_keep ), .C(\notGate[400]_keep ), 
         .D(\notGate[400]_keep ), .Z(\notGate[401] )) /* synthesis syn_instantiated=1, lut_function=((!D !C !B !A)+(!D !C !B A)+(!D !C B !A)+(!D !C B A)+(!D C !B !A)+(!D C !B A)+(!D C B !A)+(!D C B A)), LSE_LINE_FILE_ID=3, LSE_LCOL=13, LSE_RCOL=44, LSE_LLINE=32, LSE_RLINE=32 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(11[2:53])
    defparam I1.init = 16'b0000000011111111;
    
endmodule
//
// Verilog Description of module inverter_U664
//

module inverter_U664 (\notGate[399]_keep , \notGate[400] ) /* synthesis syn_module_defined=1 */ ;
    input \notGate[399]_keep ;
    output \notGate[400] ;
    
    wire \notGate[399]_keep  /* synthesis alspreserve=1 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(25[15:22])
    
    LUT4 I1 (.A(\notGate[399]_keep ), .B(\notGate[399]_keep ), .C(\notGate[399]_keep ), 
         .D(\notGate[399]_keep ), .Z(\notGate[400] )) /* synthesis syn_instantiated=1, lut_function=((!D !C !B !A)+(!D !C !B A)+(!D !C B !A)+(!D !C B A)+(!D C !B !A)+(!D C !B A)+(!D C B !A)+(!D C B A)), LSE_LINE_FILE_ID=3, LSE_LCOL=13, LSE_RCOL=44, LSE_LLINE=32, LSE_RLINE=32 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(11[2:53])
    defparam I1.init = 16'b0000000011111111;
    
endmodule
//
// Verilog Description of module inverter_U665
//

module inverter_U665 (\notGate[2]_keep , \notGate[3] ) /* synthesis syn_module_defined=1 */ ;
    input \notGate[2]_keep ;
    output \notGate[3] ;
    
    wire \notGate[2]_keep  /* synthesis alspreserve=1 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(25[15:22])
    
    LUT4 I1 (.A(\notGate[2]_keep ), .B(\notGate[2]_keep ), .C(\notGate[2]_keep ), 
         .D(\notGate[2]_keep ), .Z(\notGate[3] )) /* synthesis syn_instantiated=1, lut_function=((!D !C !B !A)+(!D !C !B A)+(!D !C B !A)+(!D !C B A)+(!D C !B !A)+(!D C !B A)+(!D C B !A)+(!D C B A)), LSE_LINE_FILE_ID=3, LSE_LCOL=13, LSE_RCOL=44, LSE_LLINE=32, LSE_RLINE=32 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(11[2:53])
    defparam I1.init = 16'b0000000011111111;
    
endmodule
//
// Verilog Description of module inverter_U666
//

module inverter_U666 (\notGate[38]_keep , \notGate[39] ) /* synthesis syn_module_defined=1 */ ;
    input \notGate[38]_keep ;
    output \notGate[39] ;
    
    wire \notGate[38]_keep  /* synthesis alspreserve=1 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(25[15:22])
    
    LUT4 I1 (.A(\notGate[38]_keep ), .B(\notGate[38]_keep ), .C(\notGate[38]_keep ), 
         .D(\notGate[38]_keep ), .Z(\notGate[39] )) /* synthesis syn_instantiated=1, lut_function=((!D !C !B !A)+(!D !C !B A)+(!D !C B !A)+(!D !C B A)+(!D C !B !A)+(!D C !B A)+(!D C B !A)+(!D C B A)), LSE_LINE_FILE_ID=3, LSE_LCOL=13, LSE_RCOL=44, LSE_LLINE=32, LSE_RLINE=32 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(11[2:53])
    defparam I1.init = 16'b0000000011111111;
    
endmodule
//
// Verilog Description of module inverter_U667
//

module inverter_U667 (\notGate[398]_keep , \notGate[399] ) /* synthesis syn_module_defined=1 */ ;
    input \notGate[398]_keep ;
    output \notGate[399] ;
    
    wire \notGate[398]_keep  /* synthesis alspreserve=1 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(25[15:22])
    
    LUT4 I1 (.A(\notGate[398]_keep ), .B(\notGate[398]_keep ), .C(\notGate[398]_keep ), 
         .D(\notGate[398]_keep ), .Z(\notGate[399] )) /* synthesis syn_instantiated=1, lut_function=((!D !C !B !A)+(!D !C !B A)+(!D !C B !A)+(!D !C B A)+(!D C !B !A)+(!D C !B A)+(!D C B !A)+(!D C B A)), LSE_LINE_FILE_ID=3, LSE_LCOL=13, LSE_RCOL=44, LSE_LLINE=32, LSE_RLINE=32 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(11[2:53])
    defparam I1.init = 16'b0000000011111111;
    
endmodule
//
// Verilog Description of module inverter_U668
//

module inverter_U668 (\notGate[397]_keep , \notGate[398] ) /* synthesis syn_module_defined=1 */ ;
    input \notGate[397]_keep ;
    output \notGate[398] ;
    
    wire \notGate[397]_keep  /* synthesis alspreserve=1 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(25[15:22])
    
    LUT4 I1 (.A(\notGate[397]_keep ), .B(\notGate[397]_keep ), .C(\notGate[397]_keep ), 
         .D(\notGate[397]_keep ), .Z(\notGate[398] )) /* synthesis syn_instantiated=1, lut_function=((!D !C !B !A)+(!D !C !B A)+(!D !C B !A)+(!D !C B A)+(!D C !B !A)+(!D C !B A)+(!D C B !A)+(!D C B A)), LSE_LINE_FILE_ID=3, LSE_LCOL=13, LSE_RCOL=44, LSE_LLINE=32, LSE_RLINE=32 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(11[2:53])
    defparam I1.init = 16'b0000000011111111;
    
endmodule
//
// Verilog Description of module inverter_U669
//

module inverter_U669 (\notGate[396]_keep , \notGate[397] ) /* synthesis syn_module_defined=1 */ ;
    input \notGate[396]_keep ;
    output \notGate[397] ;
    
    wire \notGate[396]_keep  /* synthesis alspreserve=1 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(25[15:22])
    
    LUT4 I1 (.A(\notGate[396]_keep ), .B(\notGate[396]_keep ), .C(\notGate[396]_keep ), 
         .D(\notGate[396]_keep ), .Z(\notGate[397] )) /* synthesis syn_instantiated=1, lut_function=((!D !C !B !A)+(!D !C !B A)+(!D !C B !A)+(!D !C B A)+(!D C !B !A)+(!D C !B A)+(!D C B !A)+(!D C B A)), LSE_LINE_FILE_ID=3, LSE_LCOL=13, LSE_RCOL=44, LSE_LLINE=32, LSE_RLINE=32 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(11[2:53])
    defparam I1.init = 16'b0000000011111111;
    
endmodule
//
// Verilog Description of module inverter_U670
//

module inverter_U670 (\notGate[395]_keep , \notGate[396] ) /* synthesis syn_module_defined=1 */ ;
    input \notGate[395]_keep ;
    output \notGate[396] ;
    
    wire \notGate[395]_keep  /* synthesis alspreserve=1 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(25[15:22])
    
    LUT4 I1 (.A(\notGate[395]_keep ), .B(\notGate[395]_keep ), .C(\notGate[395]_keep ), 
         .D(\notGate[395]_keep ), .Z(\notGate[396] )) /* synthesis syn_instantiated=1, lut_function=((!D !C !B !A)+(!D !C !B A)+(!D !C B !A)+(!D !C B A)+(!D C !B !A)+(!D C !B A)+(!D C B !A)+(!D C B A)), LSE_LINE_FILE_ID=3, LSE_LCOL=13, LSE_RCOL=44, LSE_LLINE=32, LSE_RLINE=32 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(11[2:53])
    defparam I1.init = 16'b0000000011111111;
    
endmodule
//
// Verilog Description of module inverter_U671
//

module inverter_U671 (\notGate[394]_keep , \notGate[395] ) /* synthesis syn_module_defined=1 */ ;
    input \notGate[394]_keep ;
    output \notGate[395] ;
    
    wire \notGate[394]_keep  /* synthesis alspreserve=1 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(25[15:22])
    
    LUT4 I1 (.A(\notGate[394]_keep ), .B(\notGate[394]_keep ), .C(\notGate[394]_keep ), 
         .D(\notGate[394]_keep ), .Z(\notGate[395] )) /* synthesis syn_instantiated=1, lut_function=((!D !C !B !A)+(!D !C !B A)+(!D !C B !A)+(!D !C B A)+(!D C !B !A)+(!D C !B A)+(!D C B !A)+(!D C B A)), LSE_LINE_FILE_ID=3, LSE_LCOL=13, LSE_RCOL=44, LSE_LLINE=32, LSE_RLINE=32 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(11[2:53])
    defparam I1.init = 16'b0000000011111111;
    
endmodule
//
// Verilog Description of module inverter_U672
//

module inverter_U672 (\notGate[393]_keep , \notGate[394] ) /* synthesis syn_module_defined=1 */ ;
    input \notGate[393]_keep ;
    output \notGate[394] ;
    
    wire \notGate[393]_keep  /* synthesis alspreserve=1 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(25[15:22])
    
    LUT4 I1 (.A(\notGate[393]_keep ), .B(\notGate[393]_keep ), .C(\notGate[393]_keep ), 
         .D(\notGate[393]_keep ), .Z(\notGate[394] )) /* synthesis syn_instantiated=1, lut_function=((!D !C !B !A)+(!D !C !B A)+(!D !C B !A)+(!D !C B A)+(!D C !B !A)+(!D C !B A)+(!D C B !A)+(!D C B A)), LSE_LINE_FILE_ID=3, LSE_LCOL=13, LSE_RCOL=44, LSE_LLINE=32, LSE_RLINE=32 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(11[2:53])
    defparam I1.init = 16'b0000000011111111;
    
endmodule
//
// Verilog Description of module inverter_U673
//

module inverter_U673 (\notGate[392]_keep , \notGate[393] ) /* synthesis syn_module_defined=1 */ ;
    input \notGate[392]_keep ;
    output \notGate[393] ;
    
    wire \notGate[392]_keep  /* synthesis alspreserve=1 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(25[15:22])
    
    LUT4 I1 (.A(\notGate[392]_keep ), .B(\notGate[392]_keep ), .C(\notGate[392]_keep ), 
         .D(\notGate[392]_keep ), .Z(\notGate[393] )) /* synthesis syn_instantiated=1, lut_function=((!D !C !B !A)+(!D !C !B A)+(!D !C B !A)+(!D !C B A)+(!D C !B !A)+(!D C !B A)+(!D C B !A)+(!D C B A)), LSE_LINE_FILE_ID=3, LSE_LCOL=13, LSE_RCOL=44, LSE_LLINE=32, LSE_RLINE=32 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(11[2:53])
    defparam I1.init = 16'b0000000011111111;
    
endmodule
//
// Verilog Description of module inverter_U674
//

module inverter_U674 (\notGate[391]_keep , \notGate[392] ) /* synthesis syn_module_defined=1 */ ;
    input \notGate[391]_keep ;
    output \notGate[392] ;
    
    wire \notGate[391]_keep  /* synthesis alspreserve=1 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(25[15:22])
    
    LUT4 I1 (.A(\notGate[391]_keep ), .B(\notGate[391]_keep ), .C(\notGate[391]_keep ), 
         .D(\notGate[391]_keep ), .Z(\notGate[392] )) /* synthesis syn_instantiated=1, lut_function=((!D !C !B !A)+(!D !C !B A)+(!D !C B !A)+(!D !C B A)+(!D C !B !A)+(!D C !B A)+(!D C B !A)+(!D C B A)), LSE_LINE_FILE_ID=3, LSE_LCOL=13, LSE_RCOL=44, LSE_LLINE=32, LSE_RLINE=32 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(11[2:53])
    defparam I1.init = 16'b0000000011111111;
    
endmodule
//
// Verilog Description of module inverter_U675
//

module inverter_U675 (\notGate[390]_keep , \notGate[391] ) /* synthesis syn_module_defined=1 */ ;
    input \notGate[390]_keep ;
    output \notGate[391] ;
    
    wire \notGate[390]_keep  /* synthesis alspreserve=1 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(25[15:22])
    
    LUT4 I1 (.A(\notGate[390]_keep ), .B(\notGate[390]_keep ), .C(\notGate[390]_keep ), 
         .D(\notGate[390]_keep ), .Z(\notGate[391] )) /* synthesis syn_instantiated=1, lut_function=((!D !C !B !A)+(!D !C !B A)+(!D !C B !A)+(!D !C B A)+(!D C !B !A)+(!D C !B A)+(!D C B !A)+(!D C B A)), LSE_LINE_FILE_ID=3, LSE_LCOL=13, LSE_RCOL=44, LSE_LLINE=32, LSE_RLINE=32 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(11[2:53])
    defparam I1.init = 16'b0000000011111111;
    
endmodule
//
// Verilog Description of module inverter_U676
//

module inverter_U676 (\notGate[389]_keep , \notGate[390] ) /* synthesis syn_module_defined=1 */ ;
    input \notGate[389]_keep ;
    output \notGate[390] ;
    
    wire \notGate[389]_keep  /* synthesis alspreserve=1 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(25[15:22])
    
    LUT4 I1 (.A(\notGate[389]_keep ), .B(\notGate[389]_keep ), .C(\notGate[389]_keep ), 
         .D(\notGate[389]_keep ), .Z(\notGate[390] )) /* synthesis syn_instantiated=1, lut_function=((!D !C !B !A)+(!D !C !B A)+(!D !C B !A)+(!D !C B A)+(!D C !B !A)+(!D C !B A)+(!D C B !A)+(!D C B A)), LSE_LINE_FILE_ID=3, LSE_LCOL=13, LSE_RCOL=44, LSE_LLINE=32, LSE_RLINE=32 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(11[2:53])
    defparam I1.init = 16'b0000000011111111;
    
endmodule
//
// Verilog Description of module inverter_U677
//

module inverter_U677 (\notGate[37]_keep , \notGate[38] ) /* synthesis syn_module_defined=1 */ ;
    input \notGate[37]_keep ;
    output \notGate[38] ;
    
    wire \notGate[37]_keep  /* synthesis alspreserve=1 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(25[15:22])
    
    LUT4 I1 (.A(\notGate[37]_keep ), .B(\notGate[37]_keep ), .C(\notGate[37]_keep ), 
         .D(\notGate[37]_keep ), .Z(\notGate[38] )) /* synthesis syn_instantiated=1, lut_function=((!D !C !B !A)+(!D !C !B A)+(!D !C B !A)+(!D !C B A)+(!D C !B !A)+(!D C !B A)+(!D C B !A)+(!D C B A)), LSE_LINE_FILE_ID=3, LSE_LCOL=13, LSE_RCOL=44, LSE_LLINE=32, LSE_RLINE=32 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(11[2:53])
    defparam I1.init = 16'b0000000011111111;
    
endmodule
//
// Verilog Description of module inverter_U678
//

module inverter_U678 (\notGate[388]_keep , \notGate[389] ) /* synthesis syn_module_defined=1 */ ;
    input \notGate[388]_keep ;
    output \notGate[389] ;
    
    wire \notGate[388]_keep  /* synthesis alspreserve=1 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(25[15:22])
    
    LUT4 I1 (.A(\notGate[388]_keep ), .B(\notGate[388]_keep ), .C(\notGate[388]_keep ), 
         .D(\notGate[388]_keep ), .Z(\notGate[389] )) /* synthesis syn_instantiated=1, lut_function=((!D !C !B !A)+(!D !C !B A)+(!D !C B !A)+(!D !C B A)+(!D C !B !A)+(!D C !B A)+(!D C B !A)+(!D C B A)), LSE_LINE_FILE_ID=3, LSE_LCOL=13, LSE_RCOL=44, LSE_LLINE=32, LSE_RLINE=32 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(11[2:53])
    defparam I1.init = 16'b0000000011111111;
    
endmodule
//
// Verilog Description of module inverter_U679
//

module inverter_U679 (\notGate[387]_keep , \notGate[388] ) /* synthesis syn_module_defined=1 */ ;
    input \notGate[387]_keep ;
    output \notGate[388] ;
    
    wire \notGate[387]_keep  /* synthesis alspreserve=1 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(25[15:22])
    
    LUT4 I1 (.A(\notGate[387]_keep ), .B(\notGate[387]_keep ), .C(\notGate[387]_keep ), 
         .D(\notGate[387]_keep ), .Z(\notGate[388] )) /* synthesis syn_instantiated=1, lut_function=((!D !C !B !A)+(!D !C !B A)+(!D !C B !A)+(!D !C B A)+(!D C !B !A)+(!D C !B A)+(!D C B !A)+(!D C B A)), LSE_LINE_FILE_ID=3, LSE_LCOL=13, LSE_RCOL=44, LSE_LLINE=32, LSE_RLINE=32 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(11[2:53])
    defparam I1.init = 16'b0000000011111111;
    
endmodule
//
// Verilog Description of module inverter_U680
//

module inverter_U680 (\notGate[386]_keep , \notGate[387] ) /* synthesis syn_module_defined=1 */ ;
    input \notGate[386]_keep ;
    output \notGate[387] ;
    
    wire \notGate[386]_keep  /* synthesis alspreserve=1 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(25[15:22])
    
    LUT4 I1 (.A(\notGate[386]_keep ), .B(\notGate[386]_keep ), .C(\notGate[386]_keep ), 
         .D(\notGate[386]_keep ), .Z(\notGate[387] )) /* synthesis syn_instantiated=1, lut_function=((!D !C !B !A)+(!D !C !B A)+(!D !C B !A)+(!D !C B A)+(!D C !B !A)+(!D C !B A)+(!D C B !A)+(!D C B A)), LSE_LINE_FILE_ID=3, LSE_LCOL=13, LSE_RCOL=44, LSE_LLINE=32, LSE_RLINE=32 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(11[2:53])
    defparam I1.init = 16'b0000000011111111;
    
endmodule
//
// Verilog Description of module inverter_U681
//

module inverter_U681 (\notGate[385]_keep , \notGate[386] ) /* synthesis syn_module_defined=1 */ ;
    input \notGate[385]_keep ;
    output \notGate[386] ;
    
    wire \notGate[385]_keep  /* synthesis alspreserve=1 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(25[15:22])
    
    LUT4 I1 (.A(\notGate[385]_keep ), .B(\notGate[385]_keep ), .C(\notGate[385]_keep ), 
         .D(\notGate[385]_keep ), .Z(\notGate[386] )) /* synthesis syn_instantiated=1, lut_function=((!D !C !B !A)+(!D !C !B A)+(!D !C B !A)+(!D !C B A)+(!D C !B !A)+(!D C !B A)+(!D C B !A)+(!D C B A)), LSE_LINE_FILE_ID=3, LSE_LCOL=13, LSE_RCOL=44, LSE_LLINE=32, LSE_RLINE=32 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(11[2:53])
    defparam I1.init = 16'b0000000011111111;
    
endmodule
//
// Verilog Description of module inverter_U682
//

module inverter_U682 (\notGate[384]_keep , \notGate[385] ) /* synthesis syn_module_defined=1 */ ;
    input \notGate[384]_keep ;
    output \notGate[385] ;
    
    wire \notGate[384]_keep  /* synthesis alspreserve=1 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(25[15:22])
    
    LUT4 I1 (.A(\notGate[384]_keep ), .B(\notGate[384]_keep ), .C(\notGate[384]_keep ), 
         .D(\notGate[384]_keep ), .Z(\notGate[385] )) /* synthesis syn_instantiated=1, lut_function=((!D !C !B !A)+(!D !C !B A)+(!D !C B !A)+(!D !C B A)+(!D C !B !A)+(!D C !B A)+(!D C B !A)+(!D C B A)), LSE_LINE_FILE_ID=3, LSE_LCOL=13, LSE_RCOL=44, LSE_LLINE=32, LSE_RLINE=32 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(11[2:53])
    defparam I1.init = 16'b0000000011111111;
    
endmodule
//
// Verilog Description of module inverter_U683
//

module inverter_U683 (\notGate[383]_keep , \notGate[384] ) /* synthesis syn_module_defined=1 */ ;
    input \notGate[383]_keep ;
    output \notGate[384] ;
    
    wire \notGate[383]_keep  /* synthesis alspreserve=1 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(25[15:22])
    
    LUT4 I1 (.A(\notGate[383]_keep ), .B(\notGate[383]_keep ), .C(\notGate[383]_keep ), 
         .D(\notGate[383]_keep ), .Z(\notGate[384] )) /* synthesis syn_instantiated=1, lut_function=((!D !C !B !A)+(!D !C !B A)+(!D !C B !A)+(!D !C B A)+(!D C !B !A)+(!D C !B A)+(!D C B !A)+(!D C B A)), LSE_LINE_FILE_ID=3, LSE_LCOL=13, LSE_RCOL=44, LSE_LLINE=32, LSE_RLINE=32 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(11[2:53])
    defparam I1.init = 16'b0000000011111111;
    
endmodule
//
// Verilog Description of module inverter_U684
//

module inverter_U684 (\notGate[382]_keep , \notGate[383] ) /* synthesis syn_module_defined=1 */ ;
    input \notGate[382]_keep ;
    output \notGate[383] ;
    
    wire \notGate[382]_keep  /* synthesis alspreserve=1 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(25[15:22])
    
    LUT4 I1 (.A(\notGate[382]_keep ), .B(\notGate[382]_keep ), .C(\notGate[382]_keep ), 
         .D(\notGate[382]_keep ), .Z(\notGate[383] )) /* synthesis syn_instantiated=1, lut_function=((!D !C !B !A)+(!D !C !B A)+(!D !C B !A)+(!D !C B A)+(!D C !B !A)+(!D C !B A)+(!D C B !A)+(!D C B A)), LSE_LINE_FILE_ID=3, LSE_LCOL=13, LSE_RCOL=44, LSE_LLINE=32, LSE_RLINE=32 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(11[2:53])
    defparam I1.init = 16'b0000000011111111;
    
endmodule
//
// Verilog Description of module inverter_U685
//

module inverter_U685 (\notGate[381]_keep , \notGate[382] ) /* synthesis syn_module_defined=1 */ ;
    input \notGate[381]_keep ;
    output \notGate[382] ;
    
    wire \notGate[381]_keep  /* synthesis alspreserve=1 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(25[15:22])
    
    LUT4 I1 (.A(\notGate[381]_keep ), .B(\notGate[381]_keep ), .C(\notGate[381]_keep ), 
         .D(\notGate[381]_keep ), .Z(\notGate[382] )) /* synthesis syn_instantiated=1, lut_function=((!D !C !B !A)+(!D !C !B A)+(!D !C B !A)+(!D !C B A)+(!D C !B !A)+(!D C !B A)+(!D C B !A)+(!D C B A)), LSE_LINE_FILE_ID=3, LSE_LCOL=13, LSE_RCOL=44, LSE_LLINE=32, LSE_RLINE=32 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(11[2:53])
    defparam I1.init = 16'b0000000011111111;
    
endmodule
//
// Verilog Description of module inverter_U686
//

module inverter_U686 (\notGate[380]_keep , \notGate[381] ) /* synthesis syn_module_defined=1 */ ;
    input \notGate[380]_keep ;
    output \notGate[381] ;
    
    wire \notGate[380]_keep  /* synthesis alspreserve=1 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(25[15:22])
    
    LUT4 I1 (.A(\notGate[380]_keep ), .B(\notGate[380]_keep ), .C(\notGate[380]_keep ), 
         .D(\notGate[380]_keep ), .Z(\notGate[381] )) /* synthesis syn_instantiated=1, lut_function=((!D !C !B !A)+(!D !C !B A)+(!D !C B !A)+(!D !C B A)+(!D C !B !A)+(!D C !B A)+(!D C B !A)+(!D C B A)), LSE_LINE_FILE_ID=3, LSE_LCOL=13, LSE_RCOL=44, LSE_LLINE=32, LSE_RLINE=32 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(11[2:53])
    defparam I1.init = 16'b0000000011111111;
    
endmodule
//
// Verilog Description of module inverter_U687
//

module inverter_U687 (\notGate[379]_keep , \notGate[380] ) /* synthesis syn_module_defined=1 */ ;
    input \notGate[379]_keep ;
    output \notGate[380] ;
    
    wire \notGate[379]_keep  /* synthesis alspreserve=1 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(25[15:22])
    
    LUT4 I1 (.A(\notGate[379]_keep ), .B(\notGate[379]_keep ), .C(\notGate[379]_keep ), 
         .D(\notGate[379]_keep ), .Z(\notGate[380] )) /* synthesis syn_instantiated=1, lut_function=((!D !C !B !A)+(!D !C !B A)+(!D !C B !A)+(!D !C B A)+(!D C !B !A)+(!D C !B A)+(!D C B !A)+(!D C B A)), LSE_LINE_FILE_ID=3, LSE_LCOL=13, LSE_RCOL=44, LSE_LLINE=32, LSE_RLINE=32 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(11[2:53])
    defparam I1.init = 16'b0000000011111111;
    
endmodule
//
// Verilog Description of module inverter_U688
//

module inverter_U688 (\notGate[36]_keep , \notGate[37] ) /* synthesis syn_module_defined=1 */ ;
    input \notGate[36]_keep ;
    output \notGate[37] ;
    
    wire \notGate[36]_keep  /* synthesis alspreserve=1 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(25[15:22])
    
    LUT4 I1 (.A(\notGate[36]_keep ), .B(\notGate[36]_keep ), .C(\notGate[36]_keep ), 
         .D(\notGate[36]_keep ), .Z(\notGate[37] )) /* synthesis syn_instantiated=1, lut_function=((!D !C !B !A)+(!D !C !B A)+(!D !C B !A)+(!D !C B A)+(!D C !B !A)+(!D C !B A)+(!D C B !A)+(!D C B A)), LSE_LINE_FILE_ID=3, LSE_LCOL=13, LSE_RCOL=44, LSE_LLINE=32, LSE_RLINE=32 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(11[2:53])
    defparam I1.init = 16'b0000000011111111;
    
endmodule
//
// Verilog Description of module inverter_U689
//

module inverter_U689 (\notGate[378]_keep , \notGate[379] ) /* synthesis syn_module_defined=1 */ ;
    input \notGate[378]_keep ;
    output \notGate[379] ;
    
    wire \notGate[378]_keep  /* synthesis alspreserve=1 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(25[15:22])
    
    LUT4 I1 (.A(\notGate[378]_keep ), .B(\notGate[378]_keep ), .C(\notGate[378]_keep ), 
         .D(\notGate[378]_keep ), .Z(\notGate[379] )) /* synthesis syn_instantiated=1, lut_function=((!D !C !B !A)+(!D !C !B A)+(!D !C B !A)+(!D !C B A)+(!D C !B !A)+(!D C !B A)+(!D C B !A)+(!D C B A)), LSE_LINE_FILE_ID=3, LSE_LCOL=13, LSE_RCOL=44, LSE_LLINE=32, LSE_RLINE=32 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(11[2:53])
    defparam I1.init = 16'b0000000011111111;
    
endmodule
//
// Verilog Description of module inverter_U690
//

module inverter_U690 (\notGate[377]_keep , \notGate[378] ) /* synthesis syn_module_defined=1 */ ;
    input \notGate[377]_keep ;
    output \notGate[378] ;
    
    wire \notGate[377]_keep  /* synthesis alspreserve=1 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(25[15:22])
    
    LUT4 I1 (.A(\notGate[377]_keep ), .B(\notGate[377]_keep ), .C(\notGate[377]_keep ), 
         .D(\notGate[377]_keep ), .Z(\notGate[378] )) /* synthesis syn_instantiated=1, lut_function=((!D !C !B !A)+(!D !C !B A)+(!D !C B !A)+(!D !C B A)+(!D C !B !A)+(!D C !B A)+(!D C B !A)+(!D C B A)), LSE_LINE_FILE_ID=3, LSE_LCOL=13, LSE_RCOL=44, LSE_LLINE=32, LSE_RLINE=32 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(11[2:53])
    defparam I1.init = 16'b0000000011111111;
    
endmodule
//
// Verilog Description of module inverter_U691
//

module inverter_U691 (\notGate[376]_keep , \notGate[377] ) /* synthesis syn_module_defined=1 */ ;
    input \notGate[376]_keep ;
    output \notGate[377] ;
    
    wire \notGate[376]_keep  /* synthesis alspreserve=1 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(25[15:22])
    
    LUT4 I1 (.A(\notGate[376]_keep ), .B(\notGate[376]_keep ), .C(\notGate[376]_keep ), 
         .D(\notGate[376]_keep ), .Z(\notGate[377] )) /* synthesis syn_instantiated=1, lut_function=((!D !C !B !A)+(!D !C !B A)+(!D !C B !A)+(!D !C B A)+(!D C !B !A)+(!D C !B A)+(!D C B !A)+(!D C B A)), LSE_LINE_FILE_ID=3, LSE_LCOL=13, LSE_RCOL=44, LSE_LLINE=32, LSE_RLINE=32 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(11[2:53])
    defparam I1.init = 16'b0000000011111111;
    
endmodule
//
// Verilog Description of module inverter_U692
//

module inverter_U692 (\notGate[375]_keep , \notGate[376] ) /* synthesis syn_module_defined=1 */ ;
    input \notGate[375]_keep ;
    output \notGate[376] ;
    
    wire \notGate[375]_keep  /* synthesis alspreserve=1 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(25[15:22])
    
    LUT4 I1 (.A(\notGate[375]_keep ), .B(\notGate[375]_keep ), .C(\notGate[375]_keep ), 
         .D(\notGate[375]_keep ), .Z(\notGate[376] )) /* synthesis syn_instantiated=1, lut_function=((!D !C !B !A)+(!D !C !B A)+(!D !C B !A)+(!D !C B A)+(!D C !B !A)+(!D C !B A)+(!D C B !A)+(!D C B A)), LSE_LINE_FILE_ID=3, LSE_LCOL=13, LSE_RCOL=44, LSE_LLINE=32, LSE_RLINE=32 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(11[2:53])
    defparam I1.init = 16'b0000000011111111;
    
endmodule
//
// Verilog Description of module inverter_U693
//

module inverter_U693 (\notGate[374]_keep , \notGate[375] ) /* synthesis syn_module_defined=1 */ ;
    input \notGate[374]_keep ;
    output \notGate[375] ;
    
    wire \notGate[374]_keep  /* synthesis alspreserve=1 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(25[15:22])
    
    LUT4 I1 (.A(\notGate[374]_keep ), .B(\notGate[374]_keep ), .C(\notGate[374]_keep ), 
         .D(\notGate[374]_keep ), .Z(\notGate[375] )) /* synthesis syn_instantiated=1, lut_function=((!D !C !B !A)+(!D !C !B A)+(!D !C B !A)+(!D !C B A)+(!D C !B !A)+(!D C !B A)+(!D C B !A)+(!D C B A)), LSE_LINE_FILE_ID=3, LSE_LCOL=13, LSE_RCOL=44, LSE_LLINE=32, LSE_RLINE=32 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(11[2:53])
    defparam I1.init = 16'b0000000011111111;
    
endmodule
//
// Verilog Description of module inverter_U694
//

module inverter_U694 (\notGate[373]_keep , \notGate[374] ) /* synthesis syn_module_defined=1 */ ;
    input \notGate[373]_keep ;
    output \notGate[374] ;
    
    wire \notGate[373]_keep  /* synthesis alspreserve=1 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(25[15:22])
    
    LUT4 I1 (.A(\notGate[373]_keep ), .B(\notGate[373]_keep ), .C(\notGate[373]_keep ), 
         .D(\notGate[373]_keep ), .Z(\notGate[374] )) /* synthesis syn_instantiated=1, lut_function=((!D !C !B !A)+(!D !C !B A)+(!D !C B !A)+(!D !C B A)+(!D C !B !A)+(!D C !B A)+(!D C B !A)+(!D C B A)), LSE_LINE_FILE_ID=3, LSE_LCOL=13, LSE_RCOL=44, LSE_LLINE=32, LSE_RLINE=32 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(11[2:53])
    defparam I1.init = 16'b0000000011111111;
    
endmodule
//
// Verilog Description of module inverter_U695
//

module inverter_U695 (\notGate[372]_keep , \notGate[373] ) /* synthesis syn_module_defined=1 */ ;
    input \notGate[372]_keep ;
    output \notGate[373] ;
    
    wire \notGate[372]_keep  /* synthesis alspreserve=1 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(25[15:22])
    
    LUT4 I1 (.A(\notGate[372]_keep ), .B(\notGate[372]_keep ), .C(\notGate[372]_keep ), 
         .D(\notGate[372]_keep ), .Z(\notGate[373] )) /* synthesis syn_instantiated=1, lut_function=((!D !C !B !A)+(!D !C !B A)+(!D !C B !A)+(!D !C B A)+(!D C !B !A)+(!D C !B A)+(!D C B !A)+(!D C B A)), LSE_LINE_FILE_ID=3, LSE_LCOL=13, LSE_RCOL=44, LSE_LLINE=32, LSE_RLINE=32 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(11[2:53])
    defparam I1.init = 16'b0000000011111111;
    
endmodule
//
// Verilog Description of module inverter_U696
//

module inverter_U696 (\notGate[371]_keep , \notGate[372] ) /* synthesis syn_module_defined=1 */ ;
    input \notGate[371]_keep ;
    output \notGate[372] ;
    
    wire \notGate[371]_keep  /* synthesis alspreserve=1 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(25[15:22])
    
    LUT4 I1 (.A(\notGate[371]_keep ), .B(\notGate[371]_keep ), .C(\notGate[371]_keep ), 
         .D(\notGate[371]_keep ), .Z(\notGate[372] )) /* synthesis syn_instantiated=1, lut_function=((!D !C !B !A)+(!D !C !B A)+(!D !C B !A)+(!D !C B A)+(!D C !B !A)+(!D C !B A)+(!D C B !A)+(!D C B A)), LSE_LINE_FILE_ID=3, LSE_LCOL=13, LSE_RCOL=44, LSE_LLINE=32, LSE_RLINE=32 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(11[2:53])
    defparam I1.init = 16'b0000000011111111;
    
endmodule
//
// Verilog Description of module inverter_U697
//

module inverter_U697 (\notGate[370]_keep , \notGate[371] ) /* synthesis syn_module_defined=1 */ ;
    input \notGate[370]_keep ;
    output \notGate[371] ;
    
    wire \notGate[370]_keep  /* synthesis alspreserve=1 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(25[15:22])
    
    LUT4 I1 (.A(\notGate[370]_keep ), .B(\notGate[370]_keep ), .C(\notGate[370]_keep ), 
         .D(\notGate[370]_keep ), .Z(\notGate[371] )) /* synthesis syn_instantiated=1, lut_function=((!D !C !B !A)+(!D !C !B A)+(!D !C B !A)+(!D !C B A)+(!D C !B !A)+(!D C !B A)+(!D C B !A)+(!D C B A)), LSE_LINE_FILE_ID=3, LSE_LCOL=13, LSE_RCOL=44, LSE_LLINE=32, LSE_RLINE=32 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(11[2:53])
    defparam I1.init = 16'b0000000011111111;
    
endmodule
//
// Verilog Description of module inverter_U698
//

module inverter_U698 (\notGate[369]_keep , \notGate[370] ) /* synthesis syn_module_defined=1 */ ;
    input \notGate[369]_keep ;
    output \notGate[370] ;
    
    wire \notGate[369]_keep  /* synthesis alspreserve=1 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(25[15:22])
    
    LUT4 I1 (.A(\notGate[369]_keep ), .B(\notGate[369]_keep ), .C(\notGate[369]_keep ), 
         .D(\notGate[369]_keep ), .Z(\notGate[370] )) /* synthesis syn_instantiated=1, lut_function=((!D !C !B !A)+(!D !C !B A)+(!D !C B !A)+(!D !C B A)+(!D C !B !A)+(!D C !B A)+(!D C B !A)+(!D C B A)), LSE_LINE_FILE_ID=3, LSE_LCOL=13, LSE_RCOL=44, LSE_LLINE=32, LSE_RLINE=32 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(11[2:53])
    defparam I1.init = 16'b0000000011111111;
    
endmodule
//
// Verilog Description of module inverter_U699
//

module inverter_U699 (\notGate[35]_keep , \notGate[36] ) /* synthesis syn_module_defined=1 */ ;
    input \notGate[35]_keep ;
    output \notGate[36] ;
    
    wire \notGate[35]_keep  /* synthesis alspreserve=1 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(25[15:22])
    
    LUT4 I1 (.A(\notGate[35]_keep ), .B(\notGate[35]_keep ), .C(\notGate[35]_keep ), 
         .D(\notGate[35]_keep ), .Z(\notGate[36] )) /* synthesis syn_instantiated=1, lut_function=((!D !C !B !A)+(!D !C !B A)+(!D !C B !A)+(!D !C B A)+(!D C !B !A)+(!D C !B A)+(!D C B !A)+(!D C B A)), LSE_LINE_FILE_ID=3, LSE_LCOL=13, LSE_RCOL=44, LSE_LLINE=32, LSE_RLINE=32 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(11[2:53])
    defparam I1.init = 16'b0000000011111111;
    
endmodule
//
// Verilog Description of module inverter_U700
//

module inverter_U700 (\notGate[368]_keep , \notGate[369] ) /* synthesis syn_module_defined=1 */ ;
    input \notGate[368]_keep ;
    output \notGate[369] ;
    
    wire \notGate[368]_keep  /* synthesis alspreserve=1 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(25[15:22])
    
    LUT4 I1 (.A(\notGate[368]_keep ), .B(\notGate[368]_keep ), .C(\notGate[368]_keep ), 
         .D(\notGate[368]_keep ), .Z(\notGate[369] )) /* synthesis syn_instantiated=1, lut_function=((!D !C !B !A)+(!D !C !B A)+(!D !C B !A)+(!D !C B A)+(!D C !B !A)+(!D C !B A)+(!D C B !A)+(!D C B A)), LSE_LINE_FILE_ID=3, LSE_LCOL=13, LSE_RCOL=44, LSE_LLINE=32, LSE_RLINE=32 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(11[2:53])
    defparam I1.init = 16'b0000000011111111;
    
endmodule
//
// Verilog Description of module inverter_U701
//

module inverter_U701 (\notGate[367]_keep , \notGate[368] ) /* synthesis syn_module_defined=1 */ ;
    input \notGate[367]_keep ;
    output \notGate[368] ;
    
    wire \notGate[367]_keep  /* synthesis alspreserve=1 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(25[15:22])
    
    LUT4 I1 (.A(\notGate[367]_keep ), .B(\notGate[367]_keep ), .C(\notGate[367]_keep ), 
         .D(\notGate[367]_keep ), .Z(\notGate[368] )) /* synthesis syn_instantiated=1, lut_function=((!D !C !B !A)+(!D !C !B A)+(!D !C B !A)+(!D !C B A)+(!D C !B !A)+(!D C !B A)+(!D C B !A)+(!D C B A)), LSE_LINE_FILE_ID=3, LSE_LCOL=13, LSE_RCOL=44, LSE_LLINE=32, LSE_RLINE=32 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(11[2:53])
    defparam I1.init = 16'b0000000011111111;
    
endmodule
//
// Verilog Description of module inverter_U702
//

module inverter_U702 (\notGate[366]_keep , \notGate[367] ) /* synthesis syn_module_defined=1 */ ;
    input \notGate[366]_keep ;
    output \notGate[367] ;
    
    wire \notGate[366]_keep  /* synthesis alspreserve=1 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(25[15:22])
    
    LUT4 I1 (.A(\notGate[366]_keep ), .B(\notGate[366]_keep ), .C(\notGate[366]_keep ), 
         .D(\notGate[366]_keep ), .Z(\notGate[367] )) /* synthesis syn_instantiated=1, lut_function=((!D !C !B !A)+(!D !C !B A)+(!D !C B !A)+(!D !C B A)+(!D C !B !A)+(!D C !B A)+(!D C B !A)+(!D C B A)), LSE_LINE_FILE_ID=3, LSE_LCOL=13, LSE_RCOL=44, LSE_LLINE=32, LSE_RLINE=32 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(11[2:53])
    defparam I1.init = 16'b0000000011111111;
    
endmodule
//
// Verilog Description of module inverter_U703
//

module inverter_U703 (\notGate[365]_keep , \notGate[366] ) /* synthesis syn_module_defined=1 */ ;
    input \notGate[365]_keep ;
    output \notGate[366] ;
    
    wire \notGate[365]_keep  /* synthesis alspreserve=1 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(25[15:22])
    
    LUT4 I1 (.A(\notGate[365]_keep ), .B(\notGate[365]_keep ), .C(\notGate[365]_keep ), 
         .D(\notGate[365]_keep ), .Z(\notGate[366] )) /* synthesis syn_instantiated=1, lut_function=((!D !C !B !A)+(!D !C !B A)+(!D !C B !A)+(!D !C B A)+(!D C !B !A)+(!D C !B A)+(!D C B !A)+(!D C B A)), LSE_LINE_FILE_ID=3, LSE_LCOL=13, LSE_RCOL=44, LSE_LLINE=32, LSE_RLINE=32 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(11[2:53])
    defparam I1.init = 16'b0000000011111111;
    
endmodule
//
// Verilog Description of module inverter_U704
//

module inverter_U704 (\notGate[364]_keep , \notGate[365] ) /* synthesis syn_module_defined=1 */ ;
    input \notGate[364]_keep ;
    output \notGate[365] ;
    
    wire \notGate[364]_keep  /* synthesis alspreserve=1 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(25[15:22])
    
    LUT4 I1 (.A(\notGate[364]_keep ), .B(\notGate[364]_keep ), .C(\notGate[364]_keep ), 
         .D(\notGate[364]_keep ), .Z(\notGate[365] )) /* synthesis syn_instantiated=1, lut_function=((!D !C !B !A)+(!D !C !B A)+(!D !C B !A)+(!D !C B A)+(!D C !B !A)+(!D C !B A)+(!D C B !A)+(!D C B A)), LSE_LINE_FILE_ID=3, LSE_LCOL=13, LSE_RCOL=44, LSE_LLINE=32, LSE_RLINE=32 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(11[2:53])
    defparam I1.init = 16'b0000000011111111;
    
endmodule
//
// Verilog Description of module inverter_U705
//

module inverter_U705 (\notGate[363]_keep , \notGate[364] ) /* synthesis syn_module_defined=1 */ ;
    input \notGate[363]_keep ;
    output \notGate[364] ;
    
    wire \notGate[363]_keep  /* synthesis alspreserve=1 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(25[15:22])
    
    LUT4 I1 (.A(\notGate[363]_keep ), .B(\notGate[363]_keep ), .C(\notGate[363]_keep ), 
         .D(\notGate[363]_keep ), .Z(\notGate[364] )) /* synthesis syn_instantiated=1, lut_function=((!D !C !B !A)+(!D !C !B A)+(!D !C B !A)+(!D !C B A)+(!D C !B !A)+(!D C !B A)+(!D C B !A)+(!D C B A)), LSE_LINE_FILE_ID=3, LSE_LCOL=13, LSE_RCOL=44, LSE_LLINE=32, LSE_RLINE=32 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(11[2:53])
    defparam I1.init = 16'b0000000011111111;
    
endmodule
//
// Verilog Description of module inverter_U706
//

module inverter_U706 (\notGate[362]_keep , \notGate[363] ) /* synthesis syn_module_defined=1 */ ;
    input \notGate[362]_keep ;
    output \notGate[363] ;
    
    wire \notGate[362]_keep  /* synthesis alspreserve=1 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(25[15:22])
    
    LUT4 I1 (.A(\notGate[362]_keep ), .B(\notGate[362]_keep ), .C(\notGate[362]_keep ), 
         .D(\notGate[362]_keep ), .Z(\notGate[363] )) /* synthesis syn_instantiated=1, lut_function=((!D !C !B !A)+(!D !C !B A)+(!D !C B !A)+(!D !C B A)+(!D C !B !A)+(!D C !B A)+(!D C B !A)+(!D C B A)), LSE_LINE_FILE_ID=3, LSE_LCOL=13, LSE_RCOL=44, LSE_LLINE=32, LSE_RLINE=32 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(11[2:53])
    defparam I1.init = 16'b0000000011111111;
    
endmodule
//
// Verilog Description of module inverter_U707
//

module inverter_U707 (\notGate[361]_keep , \notGate[362] ) /* synthesis syn_module_defined=1 */ ;
    input \notGate[361]_keep ;
    output \notGate[362] ;
    
    wire \notGate[361]_keep  /* synthesis alspreserve=1 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(25[15:22])
    
    LUT4 I1 (.A(\notGate[361]_keep ), .B(\notGate[361]_keep ), .C(\notGate[361]_keep ), 
         .D(\notGate[361]_keep ), .Z(\notGate[362] )) /* synthesis syn_instantiated=1, lut_function=((!D !C !B !A)+(!D !C !B A)+(!D !C B !A)+(!D !C B A)+(!D C !B !A)+(!D C !B A)+(!D C B !A)+(!D C B A)), LSE_LINE_FILE_ID=3, LSE_LCOL=13, LSE_RCOL=44, LSE_LLINE=32, LSE_RLINE=32 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(11[2:53])
    defparam I1.init = 16'b0000000011111111;
    
endmodule
//
// Verilog Description of module inverter_U708
//

module inverter_U708 (\notGate[360]_keep , \notGate[361] ) /* synthesis syn_module_defined=1 */ ;
    input \notGate[360]_keep ;
    output \notGate[361] ;
    
    wire \notGate[360]_keep  /* synthesis alspreserve=1 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(25[15:22])
    
    LUT4 I1 (.A(\notGate[360]_keep ), .B(\notGate[360]_keep ), .C(\notGate[360]_keep ), 
         .D(\notGate[360]_keep ), .Z(\notGate[361] )) /* synthesis syn_instantiated=1, lut_function=((!D !C !B !A)+(!D !C !B A)+(!D !C B !A)+(!D !C B A)+(!D C !B !A)+(!D C !B A)+(!D C B !A)+(!D C B A)), LSE_LINE_FILE_ID=3, LSE_LCOL=13, LSE_RCOL=44, LSE_LLINE=32, LSE_RLINE=32 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(11[2:53])
    defparam I1.init = 16'b0000000011111111;
    
endmodule
//
// Verilog Description of module inverter_U709
//

module inverter_U709 (\notGate[359]_keep , \notGate[360] ) /* synthesis syn_module_defined=1 */ ;
    input \notGate[359]_keep ;
    output \notGate[360] ;
    
    wire \notGate[359]_keep  /* synthesis alspreserve=1 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(25[15:22])
    
    LUT4 I1 (.A(\notGate[359]_keep ), .B(\notGate[359]_keep ), .C(\notGate[359]_keep ), 
         .D(\notGate[359]_keep ), .Z(\notGate[360] )) /* synthesis syn_instantiated=1, lut_function=((!D !C !B !A)+(!D !C !B A)+(!D !C B !A)+(!D !C B A)+(!D C !B !A)+(!D C !B A)+(!D C B !A)+(!D C B A)), LSE_LINE_FILE_ID=3, LSE_LCOL=13, LSE_RCOL=44, LSE_LLINE=32, LSE_RLINE=32 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(11[2:53])
    defparam I1.init = 16'b0000000011111111;
    
endmodule
//
// Verilog Description of module inverter_U710
//

module inverter_U710 (\notGate[34]_keep , \notGate[35] ) /* synthesis syn_module_defined=1 */ ;
    input \notGate[34]_keep ;
    output \notGate[35] ;
    
    wire \notGate[34]_keep  /* synthesis alspreserve=1 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(25[15:22])
    
    LUT4 I1 (.A(\notGate[34]_keep ), .B(\notGate[34]_keep ), .C(\notGate[34]_keep ), 
         .D(\notGate[34]_keep ), .Z(\notGate[35] )) /* synthesis syn_instantiated=1, lut_function=((!D !C !B !A)+(!D !C !B A)+(!D !C B !A)+(!D !C B A)+(!D C !B !A)+(!D C !B A)+(!D C B !A)+(!D C B A)), LSE_LINE_FILE_ID=3, LSE_LCOL=13, LSE_RCOL=44, LSE_LLINE=32, LSE_RLINE=32 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(11[2:53])
    defparam I1.init = 16'b0000000011111111;
    
endmodule
//
// Verilog Description of module inverter_U711
//

module inverter_U711 (\notGate[358]_keep , \notGate[359] ) /* synthesis syn_module_defined=1 */ ;
    input \notGate[358]_keep ;
    output \notGate[359] ;
    
    wire \notGate[358]_keep  /* synthesis alspreserve=1 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(25[15:22])
    
    LUT4 I1 (.A(\notGate[358]_keep ), .B(\notGate[358]_keep ), .C(\notGate[358]_keep ), 
         .D(\notGate[358]_keep ), .Z(\notGate[359] )) /* synthesis syn_instantiated=1, lut_function=((!D !C !B !A)+(!D !C !B A)+(!D !C B !A)+(!D !C B A)+(!D C !B !A)+(!D C !B A)+(!D C B !A)+(!D C B A)), LSE_LINE_FILE_ID=3, LSE_LCOL=13, LSE_RCOL=44, LSE_LLINE=32, LSE_RLINE=32 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(11[2:53])
    defparam I1.init = 16'b0000000011111111;
    
endmodule
//
// Verilog Description of module inverter_U712
//

module inverter_U712 (\notGate[357]_keep , \notGate[358] ) /* synthesis syn_module_defined=1 */ ;
    input \notGate[357]_keep ;
    output \notGate[358] ;
    
    wire \notGate[357]_keep  /* synthesis alspreserve=1 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(25[15:22])
    
    LUT4 I1 (.A(\notGate[357]_keep ), .B(\notGate[357]_keep ), .C(\notGate[357]_keep ), 
         .D(\notGate[357]_keep ), .Z(\notGate[358] )) /* synthesis syn_instantiated=1, lut_function=((!D !C !B !A)+(!D !C !B A)+(!D !C B !A)+(!D !C B A)+(!D C !B !A)+(!D C !B A)+(!D C B !A)+(!D C B A)), LSE_LINE_FILE_ID=3, LSE_LCOL=13, LSE_RCOL=44, LSE_LLINE=32, LSE_RLINE=32 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(11[2:53])
    defparam I1.init = 16'b0000000011111111;
    
endmodule
//
// Verilog Description of module inverter_U713
//

module inverter_U713 (\notGate[356]_keep , \notGate[357] ) /* synthesis syn_module_defined=1 */ ;
    input \notGate[356]_keep ;
    output \notGate[357] ;
    
    wire \notGate[356]_keep  /* synthesis alspreserve=1 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(25[15:22])
    
    LUT4 I1 (.A(\notGate[356]_keep ), .B(\notGate[356]_keep ), .C(\notGate[356]_keep ), 
         .D(\notGate[356]_keep ), .Z(\notGate[357] )) /* synthesis syn_instantiated=1, lut_function=((!D !C !B !A)+(!D !C !B A)+(!D !C B !A)+(!D !C B A)+(!D C !B !A)+(!D C !B A)+(!D C B !A)+(!D C B A)), LSE_LINE_FILE_ID=3, LSE_LCOL=13, LSE_RCOL=44, LSE_LLINE=32, LSE_RLINE=32 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(11[2:53])
    defparam I1.init = 16'b0000000011111111;
    
endmodule
//
// Verilog Description of module inverter_U714
//

module inverter_U714 (\notGate[355]_keep , \notGate[356] ) /* synthesis syn_module_defined=1 */ ;
    input \notGate[355]_keep ;
    output \notGate[356] ;
    
    wire \notGate[355]_keep  /* synthesis alspreserve=1 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(25[15:22])
    
    LUT4 I1 (.A(\notGate[355]_keep ), .B(\notGate[355]_keep ), .C(\notGate[355]_keep ), 
         .D(\notGate[355]_keep ), .Z(\notGate[356] )) /* synthesis syn_instantiated=1, lut_function=((!D !C !B !A)+(!D !C !B A)+(!D !C B !A)+(!D !C B A)+(!D C !B !A)+(!D C !B A)+(!D C B !A)+(!D C B A)), LSE_LINE_FILE_ID=3, LSE_LCOL=13, LSE_RCOL=44, LSE_LLINE=32, LSE_RLINE=32 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(11[2:53])
    defparam I1.init = 16'b0000000011111111;
    
endmodule
//
// Verilog Description of module inverter_U715
//

module inverter_U715 (\notGate[354]_keep , \notGate[355] ) /* synthesis syn_module_defined=1 */ ;
    input \notGate[354]_keep ;
    output \notGate[355] ;
    
    wire \notGate[354]_keep  /* synthesis alspreserve=1 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(25[15:22])
    
    LUT4 I1 (.A(\notGate[354]_keep ), .B(\notGate[354]_keep ), .C(\notGate[354]_keep ), 
         .D(\notGate[354]_keep ), .Z(\notGate[355] )) /* synthesis syn_instantiated=1, lut_function=((!D !C !B !A)+(!D !C !B A)+(!D !C B !A)+(!D !C B A)+(!D C !B !A)+(!D C !B A)+(!D C B !A)+(!D C B A)), LSE_LINE_FILE_ID=3, LSE_LCOL=13, LSE_RCOL=44, LSE_LLINE=32, LSE_RLINE=32 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(11[2:53])
    defparam I1.init = 16'b0000000011111111;
    
endmodule
//
// Verilog Description of module inverter_U716
//

module inverter_U716 (\notGate[353]_keep , \notGate[354] ) /* synthesis syn_module_defined=1 */ ;
    input \notGate[353]_keep ;
    output \notGate[354] ;
    
    wire \notGate[353]_keep  /* synthesis alspreserve=1 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(25[15:22])
    
    LUT4 I1 (.A(\notGate[353]_keep ), .B(\notGate[353]_keep ), .C(\notGate[353]_keep ), 
         .D(\notGate[353]_keep ), .Z(\notGate[354] )) /* synthesis syn_instantiated=1, lut_function=((!D !C !B !A)+(!D !C !B A)+(!D !C B !A)+(!D !C B A)+(!D C !B !A)+(!D C !B A)+(!D C B !A)+(!D C B A)), LSE_LINE_FILE_ID=3, LSE_LCOL=13, LSE_RCOL=44, LSE_LLINE=32, LSE_RLINE=32 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(11[2:53])
    defparam I1.init = 16'b0000000011111111;
    
endmodule
//
// Verilog Description of module inverter_U717
//

module inverter_U717 (\notGate[352]_keep , \notGate[353] ) /* synthesis syn_module_defined=1 */ ;
    input \notGate[352]_keep ;
    output \notGate[353] ;
    
    wire \notGate[352]_keep  /* synthesis alspreserve=1 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(25[15:22])
    
    LUT4 I1 (.A(\notGate[352]_keep ), .B(\notGate[352]_keep ), .C(\notGate[352]_keep ), 
         .D(\notGate[352]_keep ), .Z(\notGate[353] )) /* synthesis syn_instantiated=1, lut_function=((!D !C !B !A)+(!D !C !B A)+(!D !C B !A)+(!D !C B A)+(!D C !B !A)+(!D C !B A)+(!D C B !A)+(!D C B A)), LSE_LINE_FILE_ID=3, LSE_LCOL=13, LSE_RCOL=44, LSE_LLINE=32, LSE_RLINE=32 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(11[2:53])
    defparam I1.init = 16'b0000000011111111;
    
endmodule
//
// Verilog Description of module inverter_U718
//

module inverter_U718 (\notGate[351]_keep , \notGate[352] ) /* synthesis syn_module_defined=1 */ ;
    input \notGate[351]_keep ;
    output \notGate[352] ;
    
    wire \notGate[351]_keep  /* synthesis alspreserve=1 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(25[15:22])
    
    LUT4 I1 (.A(\notGate[351]_keep ), .B(\notGate[351]_keep ), .C(\notGate[351]_keep ), 
         .D(\notGate[351]_keep ), .Z(\notGate[352] )) /* synthesis syn_instantiated=1, lut_function=((!D !C !B !A)+(!D !C !B A)+(!D !C B !A)+(!D !C B A)+(!D C !B !A)+(!D C !B A)+(!D C B !A)+(!D C B A)), LSE_LINE_FILE_ID=3, LSE_LCOL=13, LSE_RCOL=44, LSE_LLINE=32, LSE_RLINE=32 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(11[2:53])
    defparam I1.init = 16'b0000000011111111;
    
endmodule
//
// Verilog Description of module inverter_U719
//

module inverter_U719 (\notGate[350]_keep , \notGate[351] ) /* synthesis syn_module_defined=1 */ ;
    input \notGate[350]_keep ;
    output \notGate[351] ;
    
    wire \notGate[350]_keep  /* synthesis alspreserve=1 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(25[15:22])
    
    LUT4 I1 (.A(\notGate[350]_keep ), .B(\notGate[350]_keep ), .C(\notGate[350]_keep ), 
         .D(\notGate[350]_keep ), .Z(\notGate[351] )) /* synthesis syn_instantiated=1, lut_function=((!D !C !B !A)+(!D !C !B A)+(!D !C B !A)+(!D !C B A)+(!D C !B !A)+(!D C !B A)+(!D C B !A)+(!D C B A)), LSE_LINE_FILE_ID=3, LSE_LCOL=13, LSE_RCOL=44, LSE_LLINE=32, LSE_RLINE=32 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(11[2:53])
    defparam I1.init = 16'b0000000011111111;
    
endmodule
//
// Verilog Description of module inverter_U720
//

module inverter_U720 (\notGate[349]_keep , \notGate[350] ) /* synthesis syn_module_defined=1 */ ;
    input \notGate[349]_keep ;
    output \notGate[350] ;
    
    wire \notGate[349]_keep  /* synthesis alspreserve=1 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(25[15:22])
    
    LUT4 I1 (.A(\notGate[349]_keep ), .B(\notGate[349]_keep ), .C(\notGate[349]_keep ), 
         .D(\notGate[349]_keep ), .Z(\notGate[350] )) /* synthesis syn_instantiated=1, lut_function=((!D !C !B !A)+(!D !C !B A)+(!D !C B !A)+(!D !C B A)+(!D C !B !A)+(!D C !B A)+(!D C B !A)+(!D C B A)), LSE_LINE_FILE_ID=3, LSE_LCOL=13, LSE_RCOL=44, LSE_LLINE=32, LSE_RLINE=32 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(11[2:53])
    defparam I1.init = 16'b0000000011111111;
    
endmodule
//
// Verilog Description of module inverter_U721
//

module inverter_U721 (\notGate[33]_keep , \notGate[34] ) /* synthesis syn_module_defined=1 */ ;
    input \notGate[33]_keep ;
    output \notGate[34] ;
    
    wire \notGate[33]_keep  /* synthesis alspreserve=1 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(25[15:22])
    
    LUT4 I1 (.A(\notGate[33]_keep ), .B(\notGate[33]_keep ), .C(\notGate[33]_keep ), 
         .D(\notGate[33]_keep ), .Z(\notGate[34] )) /* synthesis syn_instantiated=1, lut_function=((!D !C !B !A)+(!D !C !B A)+(!D !C B !A)+(!D !C B A)+(!D C !B !A)+(!D C !B A)+(!D C B !A)+(!D C B A)), LSE_LINE_FILE_ID=3, LSE_LCOL=13, LSE_RCOL=44, LSE_LLINE=32, LSE_RLINE=32 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(11[2:53])
    defparam I1.init = 16'b0000000011111111;
    
endmodule
//
// Verilog Description of module inverter_U722
//

module inverter_U722 (\notGate[348]_keep , \notGate[349] ) /* synthesis syn_module_defined=1 */ ;
    input \notGate[348]_keep ;
    output \notGate[349] ;
    
    wire \notGate[348]_keep  /* synthesis alspreserve=1 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(25[15:22])
    
    LUT4 I1 (.A(\notGate[348]_keep ), .B(\notGate[348]_keep ), .C(\notGate[348]_keep ), 
         .D(\notGate[348]_keep ), .Z(\notGate[349] )) /* synthesis syn_instantiated=1, lut_function=((!D !C !B !A)+(!D !C !B A)+(!D !C B !A)+(!D !C B A)+(!D C !B !A)+(!D C !B A)+(!D C B !A)+(!D C B A)), LSE_LINE_FILE_ID=3, LSE_LCOL=13, LSE_RCOL=44, LSE_LLINE=32, LSE_RLINE=32 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(11[2:53])
    defparam I1.init = 16'b0000000011111111;
    
endmodule
//
// Verilog Description of module inverter_U723
//

module inverter_U723 (\notGate[347]_keep , \notGate[348] ) /* synthesis syn_module_defined=1 */ ;
    input \notGate[347]_keep ;
    output \notGate[348] ;
    
    wire \notGate[347]_keep  /* synthesis alspreserve=1 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(25[15:22])
    
    LUT4 I1 (.A(\notGate[347]_keep ), .B(\notGate[347]_keep ), .C(\notGate[347]_keep ), 
         .D(\notGate[347]_keep ), .Z(\notGate[348] )) /* synthesis syn_instantiated=1, lut_function=((!D !C !B !A)+(!D !C !B A)+(!D !C B !A)+(!D !C B A)+(!D C !B !A)+(!D C !B A)+(!D C B !A)+(!D C B A)), LSE_LINE_FILE_ID=3, LSE_LCOL=13, LSE_RCOL=44, LSE_LLINE=32, LSE_RLINE=32 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(11[2:53])
    defparam I1.init = 16'b0000000011111111;
    
endmodule
//
// Verilog Description of module inverter_U724
//

module inverter_U724 (\notGate[346]_keep , \notGate[347] ) /* synthesis syn_module_defined=1 */ ;
    input \notGate[346]_keep ;
    output \notGate[347] ;
    
    wire \notGate[346]_keep  /* synthesis alspreserve=1 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(25[15:22])
    
    LUT4 I1 (.A(\notGate[346]_keep ), .B(\notGate[346]_keep ), .C(\notGate[346]_keep ), 
         .D(\notGate[346]_keep ), .Z(\notGate[347] )) /* synthesis syn_instantiated=1, lut_function=((!D !C !B !A)+(!D !C !B A)+(!D !C B !A)+(!D !C B A)+(!D C !B !A)+(!D C !B A)+(!D C B !A)+(!D C B A)), LSE_LINE_FILE_ID=3, LSE_LCOL=13, LSE_RCOL=44, LSE_LLINE=32, LSE_RLINE=32 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(11[2:53])
    defparam I1.init = 16'b0000000011111111;
    
endmodule
//
// Verilog Description of module inverter_U725
//

module inverter_U725 (\notGate[345]_keep , \notGate[346] ) /* synthesis syn_module_defined=1 */ ;
    input \notGate[345]_keep ;
    output \notGate[346] ;
    
    wire \notGate[345]_keep  /* synthesis alspreserve=1 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(25[15:22])
    
    LUT4 I1 (.A(\notGate[345]_keep ), .B(\notGate[345]_keep ), .C(\notGate[345]_keep ), 
         .D(\notGate[345]_keep ), .Z(\notGate[346] )) /* synthesis syn_instantiated=1, lut_function=((!D !C !B !A)+(!D !C !B A)+(!D !C B !A)+(!D !C B A)+(!D C !B !A)+(!D C !B A)+(!D C B !A)+(!D C B A)), LSE_LINE_FILE_ID=3, LSE_LCOL=13, LSE_RCOL=44, LSE_LLINE=32, LSE_RLINE=32 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(11[2:53])
    defparam I1.init = 16'b0000000011111111;
    
endmodule
//
// Verilog Description of module inverter_U726
//

module inverter_U726 (\notGate[344]_keep , \notGate[345] ) /* synthesis syn_module_defined=1 */ ;
    input \notGate[344]_keep ;
    output \notGate[345] ;
    
    wire \notGate[344]_keep  /* synthesis alspreserve=1 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(25[15:22])
    
    LUT4 I1 (.A(\notGate[344]_keep ), .B(\notGate[344]_keep ), .C(\notGate[344]_keep ), 
         .D(\notGate[344]_keep ), .Z(\notGate[345] )) /* synthesis syn_instantiated=1, lut_function=((!D !C !B !A)+(!D !C !B A)+(!D !C B !A)+(!D !C B A)+(!D C !B !A)+(!D C !B A)+(!D C B !A)+(!D C B A)), LSE_LINE_FILE_ID=3, LSE_LCOL=13, LSE_RCOL=44, LSE_LLINE=32, LSE_RLINE=32 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(11[2:53])
    defparam I1.init = 16'b0000000011111111;
    
endmodule
//
// Verilog Description of module inverter_U727
//

module inverter_U727 (\notGate[343]_keep , \notGate[344] ) /* synthesis syn_module_defined=1 */ ;
    input \notGate[343]_keep ;
    output \notGate[344] ;
    
    wire \notGate[343]_keep  /* synthesis alspreserve=1 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(25[15:22])
    
    LUT4 I1 (.A(\notGate[343]_keep ), .B(\notGate[343]_keep ), .C(\notGate[343]_keep ), 
         .D(\notGate[343]_keep ), .Z(\notGate[344] )) /* synthesis syn_instantiated=1, lut_function=((!D !C !B !A)+(!D !C !B A)+(!D !C B !A)+(!D !C B A)+(!D C !B !A)+(!D C !B A)+(!D C B !A)+(!D C B A)), LSE_LINE_FILE_ID=3, LSE_LCOL=13, LSE_RCOL=44, LSE_LLINE=32, LSE_RLINE=32 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(11[2:53])
    defparam I1.init = 16'b0000000011111111;
    
endmodule
//
// Verilog Description of module inverter_U728
//

module inverter_U728 (\notGate[342]_keep , \notGate[343] ) /* synthesis syn_module_defined=1 */ ;
    input \notGate[342]_keep ;
    output \notGate[343] ;
    
    wire \notGate[342]_keep  /* synthesis alspreserve=1 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(25[15:22])
    
    LUT4 I1 (.A(\notGate[342]_keep ), .B(\notGate[342]_keep ), .C(\notGate[342]_keep ), 
         .D(\notGate[342]_keep ), .Z(\notGate[343] )) /* synthesis syn_instantiated=1, lut_function=((!D !C !B !A)+(!D !C !B A)+(!D !C B !A)+(!D !C B A)+(!D C !B !A)+(!D C !B A)+(!D C B !A)+(!D C B A)), LSE_LINE_FILE_ID=3, LSE_LCOL=13, LSE_RCOL=44, LSE_LLINE=32, LSE_RLINE=32 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(11[2:53])
    defparam I1.init = 16'b0000000011111111;
    
endmodule
//
// Verilog Description of module inverter_U729
//

module inverter_U729 (\notGate[341]_keep , \notGate[342] ) /* synthesis syn_module_defined=1 */ ;
    input \notGate[341]_keep ;
    output \notGate[342] ;
    
    wire \notGate[341]_keep  /* synthesis alspreserve=1 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(25[15:22])
    
    LUT4 I1 (.A(\notGate[341]_keep ), .B(\notGate[341]_keep ), .C(\notGate[341]_keep ), 
         .D(\notGate[341]_keep ), .Z(\notGate[342] )) /* synthesis syn_instantiated=1, lut_function=((!D !C !B !A)+(!D !C !B A)+(!D !C B !A)+(!D !C B A)+(!D C !B !A)+(!D C !B A)+(!D C B !A)+(!D C B A)), LSE_LINE_FILE_ID=3, LSE_LCOL=13, LSE_RCOL=44, LSE_LLINE=32, LSE_RLINE=32 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(11[2:53])
    defparam I1.init = 16'b0000000011111111;
    
endmodule
//
// Verilog Description of module inverter_U730
//

module inverter_U730 (\notGate[340]_keep , \notGate[341] ) /* synthesis syn_module_defined=1 */ ;
    input \notGate[340]_keep ;
    output \notGate[341] ;
    
    wire \notGate[340]_keep  /* synthesis alspreserve=1 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(25[15:22])
    
    LUT4 I1 (.A(\notGate[340]_keep ), .B(\notGate[340]_keep ), .C(\notGate[340]_keep ), 
         .D(\notGate[340]_keep ), .Z(\notGate[341] )) /* synthesis syn_instantiated=1, lut_function=((!D !C !B !A)+(!D !C !B A)+(!D !C B !A)+(!D !C B A)+(!D C !B !A)+(!D C !B A)+(!D C B !A)+(!D C B A)), LSE_LINE_FILE_ID=3, LSE_LCOL=13, LSE_RCOL=44, LSE_LLINE=32, LSE_RLINE=32 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(11[2:53])
    defparam I1.init = 16'b0000000011111111;
    
endmodule
//
// Verilog Description of module inverter_U731
//

module inverter_U731 (\notGate[339]_keep , \notGate[340] ) /* synthesis syn_module_defined=1 */ ;
    input \notGate[339]_keep ;
    output \notGate[340] ;
    
    wire \notGate[339]_keep  /* synthesis alspreserve=1 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(25[15:22])
    
    LUT4 I1 (.A(\notGate[339]_keep ), .B(\notGate[339]_keep ), .C(\notGate[339]_keep ), 
         .D(\notGate[339]_keep ), .Z(\notGate[340] )) /* synthesis syn_instantiated=1, lut_function=((!D !C !B !A)+(!D !C !B A)+(!D !C B !A)+(!D !C B A)+(!D C !B !A)+(!D C !B A)+(!D C B !A)+(!D C B A)), LSE_LINE_FILE_ID=3, LSE_LCOL=13, LSE_RCOL=44, LSE_LLINE=32, LSE_RLINE=32 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(11[2:53])
    defparam I1.init = 16'b0000000011111111;
    
endmodule
//
// Verilog Description of module inverter_U732
//

module inverter_U732 (\notGate[32]_keep , \notGate[33] ) /* synthesis syn_module_defined=1 */ ;
    input \notGate[32]_keep ;
    output \notGate[33] ;
    
    wire \notGate[32]_keep  /* synthesis alspreserve=1 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(25[15:22])
    
    LUT4 I1 (.A(\notGate[32]_keep ), .B(\notGate[32]_keep ), .C(\notGate[32]_keep ), 
         .D(\notGate[32]_keep ), .Z(\notGate[33] )) /* synthesis syn_instantiated=1, lut_function=((!D !C !B !A)+(!D !C !B A)+(!D !C B !A)+(!D !C B A)+(!D C !B !A)+(!D C !B A)+(!D C B !A)+(!D C B A)), LSE_LINE_FILE_ID=3, LSE_LCOL=13, LSE_RCOL=44, LSE_LLINE=32, LSE_RLINE=32 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(11[2:53])
    defparam I1.init = 16'b0000000011111111;
    
endmodule
//
// Verilog Description of module inverter_U733
//

module inverter_U733 (\notGate[338]_keep , \notGate[339] ) /* synthesis syn_module_defined=1 */ ;
    input \notGate[338]_keep ;
    output \notGate[339] ;
    
    wire \notGate[338]_keep  /* synthesis alspreserve=1 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(25[15:22])
    
    LUT4 I1 (.A(\notGate[338]_keep ), .B(\notGate[338]_keep ), .C(\notGate[338]_keep ), 
         .D(\notGate[338]_keep ), .Z(\notGate[339] )) /* synthesis syn_instantiated=1, lut_function=((!D !C !B !A)+(!D !C !B A)+(!D !C B !A)+(!D !C B A)+(!D C !B !A)+(!D C !B A)+(!D C B !A)+(!D C B A)), LSE_LINE_FILE_ID=3, LSE_LCOL=13, LSE_RCOL=44, LSE_LLINE=32, LSE_RLINE=32 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(11[2:53])
    defparam I1.init = 16'b0000000011111111;
    
endmodule
//
// Verilog Description of module inverter_U734
//

module inverter_U734 (\notGate[337]_keep , \notGate[338] ) /* synthesis syn_module_defined=1 */ ;
    input \notGate[337]_keep ;
    output \notGate[338] ;
    
    wire \notGate[337]_keep  /* synthesis alspreserve=1 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(25[15:22])
    
    LUT4 I1 (.A(\notGate[337]_keep ), .B(\notGate[337]_keep ), .C(\notGate[337]_keep ), 
         .D(\notGate[337]_keep ), .Z(\notGate[338] )) /* synthesis syn_instantiated=1, lut_function=((!D !C !B !A)+(!D !C !B A)+(!D !C B !A)+(!D !C B A)+(!D C !B !A)+(!D C !B A)+(!D C B !A)+(!D C B A)), LSE_LINE_FILE_ID=3, LSE_LCOL=13, LSE_RCOL=44, LSE_LLINE=32, LSE_RLINE=32 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(11[2:53])
    defparam I1.init = 16'b0000000011111111;
    
endmodule
//
// Verilog Description of module inverter_U735
//

module inverter_U735 (\notGate[336]_keep , \notGate[337] ) /* synthesis syn_module_defined=1 */ ;
    input \notGate[336]_keep ;
    output \notGate[337] ;
    
    wire \notGate[336]_keep  /* synthesis alspreserve=1 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(25[15:22])
    
    LUT4 I1 (.A(\notGate[336]_keep ), .B(\notGate[336]_keep ), .C(\notGate[336]_keep ), 
         .D(\notGate[336]_keep ), .Z(\notGate[337] )) /* synthesis syn_instantiated=1, lut_function=((!D !C !B !A)+(!D !C !B A)+(!D !C B !A)+(!D !C B A)+(!D C !B !A)+(!D C !B A)+(!D C B !A)+(!D C B A)), LSE_LINE_FILE_ID=3, LSE_LCOL=13, LSE_RCOL=44, LSE_LLINE=32, LSE_RLINE=32 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(11[2:53])
    defparam I1.init = 16'b0000000011111111;
    
endmodule
//
// Verilog Description of module inverter_U736
//

module inverter_U736 (\notGate[335]_keep , \notGate[336] ) /* synthesis syn_module_defined=1 */ ;
    input \notGate[335]_keep ;
    output \notGate[336] ;
    
    wire \notGate[335]_keep  /* synthesis alspreserve=1 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(25[15:22])
    
    LUT4 I1 (.A(\notGate[335]_keep ), .B(\notGate[335]_keep ), .C(\notGate[335]_keep ), 
         .D(\notGate[335]_keep ), .Z(\notGate[336] )) /* synthesis syn_instantiated=1, lut_function=((!D !C !B !A)+(!D !C !B A)+(!D !C B !A)+(!D !C B A)+(!D C !B !A)+(!D C !B A)+(!D C B !A)+(!D C B A)), LSE_LINE_FILE_ID=3, LSE_LCOL=13, LSE_RCOL=44, LSE_LLINE=32, LSE_RLINE=32 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(11[2:53])
    defparam I1.init = 16'b0000000011111111;
    
endmodule
//
// Verilog Description of module inverter_U737
//

module inverter_U737 (\notGate[334]_keep , \notGate[335] ) /* synthesis syn_module_defined=1 */ ;
    input \notGate[334]_keep ;
    output \notGate[335] ;
    
    wire \notGate[334]_keep  /* synthesis alspreserve=1 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(25[15:22])
    
    LUT4 I1 (.A(\notGate[334]_keep ), .B(\notGate[334]_keep ), .C(\notGate[334]_keep ), 
         .D(\notGate[334]_keep ), .Z(\notGate[335] )) /* synthesis syn_instantiated=1, lut_function=((!D !C !B !A)+(!D !C !B A)+(!D !C B !A)+(!D !C B A)+(!D C !B !A)+(!D C !B A)+(!D C B !A)+(!D C B A)), LSE_LINE_FILE_ID=3, LSE_LCOL=13, LSE_RCOL=44, LSE_LLINE=32, LSE_RLINE=32 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(11[2:53])
    defparam I1.init = 16'b0000000011111111;
    
endmodule
//
// Verilog Description of module inverter_U738
//

module inverter_U738 (\notGate[333]_keep , \notGate[334] ) /* synthesis syn_module_defined=1 */ ;
    input \notGate[333]_keep ;
    output \notGate[334] ;
    
    wire \notGate[333]_keep  /* synthesis alspreserve=1 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(25[15:22])
    
    LUT4 I1 (.A(\notGate[333]_keep ), .B(\notGate[333]_keep ), .C(\notGate[333]_keep ), 
         .D(\notGate[333]_keep ), .Z(\notGate[334] )) /* synthesis syn_instantiated=1, lut_function=((!D !C !B !A)+(!D !C !B A)+(!D !C B !A)+(!D !C B A)+(!D C !B !A)+(!D C !B A)+(!D C B !A)+(!D C B A)), LSE_LINE_FILE_ID=3, LSE_LCOL=13, LSE_RCOL=44, LSE_LLINE=32, LSE_RLINE=32 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(11[2:53])
    defparam I1.init = 16'b0000000011111111;
    
endmodule
//
// Verilog Description of module inverter_U739
//

module inverter_U739 (\notGate[332]_keep , \notGate[333] ) /* synthesis syn_module_defined=1 */ ;
    input \notGate[332]_keep ;
    output \notGate[333] ;
    
    wire \notGate[332]_keep  /* synthesis alspreserve=1 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(25[15:22])
    
    LUT4 I1 (.A(\notGate[332]_keep ), .B(\notGate[332]_keep ), .C(\notGate[332]_keep ), 
         .D(\notGate[332]_keep ), .Z(\notGate[333] )) /* synthesis syn_instantiated=1, lut_function=((!D !C !B !A)+(!D !C !B A)+(!D !C B !A)+(!D !C B A)+(!D C !B !A)+(!D C !B A)+(!D C B !A)+(!D C B A)), LSE_LINE_FILE_ID=3, LSE_LCOL=13, LSE_RCOL=44, LSE_LLINE=32, LSE_RLINE=32 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(11[2:53])
    defparam I1.init = 16'b0000000011111111;
    
endmodule
//
// Verilog Description of module inverter_U740
//

module inverter_U740 (\notGate[331]_keep , \notGate[332] ) /* synthesis syn_module_defined=1 */ ;
    input \notGate[331]_keep ;
    output \notGate[332] ;
    
    wire \notGate[331]_keep  /* synthesis alspreserve=1 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(25[15:22])
    
    LUT4 I1 (.A(\notGate[331]_keep ), .B(\notGate[331]_keep ), .C(\notGate[331]_keep ), 
         .D(\notGate[331]_keep ), .Z(\notGate[332] )) /* synthesis syn_instantiated=1, lut_function=((!D !C !B !A)+(!D !C !B A)+(!D !C B !A)+(!D !C B A)+(!D C !B !A)+(!D C !B A)+(!D C B !A)+(!D C B A)), LSE_LINE_FILE_ID=3, LSE_LCOL=13, LSE_RCOL=44, LSE_LLINE=32, LSE_RLINE=32 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(11[2:53])
    defparam I1.init = 16'b0000000011111111;
    
endmodule
//
// Verilog Description of module inverter_U741
//

module inverter_U741 (\notGate[330]_keep , \notGate[331] ) /* synthesis syn_module_defined=1 */ ;
    input \notGate[330]_keep ;
    output \notGate[331] ;
    
    wire \notGate[330]_keep  /* synthesis alspreserve=1 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(25[15:22])
    
    LUT4 I1 (.A(\notGate[330]_keep ), .B(\notGate[330]_keep ), .C(\notGate[330]_keep ), 
         .D(\notGate[330]_keep ), .Z(\notGate[331] )) /* synthesis syn_instantiated=1, lut_function=((!D !C !B !A)+(!D !C !B A)+(!D !C B !A)+(!D !C B A)+(!D C !B !A)+(!D C !B A)+(!D C B !A)+(!D C B A)), LSE_LINE_FILE_ID=3, LSE_LCOL=13, LSE_RCOL=44, LSE_LLINE=32, LSE_RLINE=32 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(11[2:53])
    defparam I1.init = 16'b0000000011111111;
    
endmodule
//
// Verilog Description of module inverter_U742
//

module inverter_U742 (\notGate[329]_keep , \notGate[330] ) /* synthesis syn_module_defined=1 */ ;
    input \notGate[329]_keep ;
    output \notGate[330] ;
    
    wire \notGate[329]_keep  /* synthesis alspreserve=1 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(25[15:22])
    
    LUT4 I1 (.A(\notGate[329]_keep ), .B(\notGate[329]_keep ), .C(\notGate[329]_keep ), 
         .D(\notGate[329]_keep ), .Z(\notGate[330] )) /* synthesis syn_instantiated=1, lut_function=((!D !C !B !A)+(!D !C !B A)+(!D !C B !A)+(!D !C B A)+(!D C !B !A)+(!D C !B A)+(!D C B !A)+(!D C B A)), LSE_LINE_FILE_ID=3, LSE_LCOL=13, LSE_RCOL=44, LSE_LLINE=32, LSE_RLINE=32 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(11[2:53])
    defparam I1.init = 16'b0000000011111111;
    
endmodule
//
// Verilog Description of module inverter_U743
//

module inverter_U743 (\notGate[31]_keep , \notGate[32] ) /* synthesis syn_module_defined=1 */ ;
    input \notGate[31]_keep ;
    output \notGate[32] ;
    
    wire \notGate[31]_keep  /* synthesis alspreserve=1 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(25[15:22])
    
    LUT4 I1 (.A(\notGate[31]_keep ), .B(\notGate[31]_keep ), .C(\notGate[31]_keep ), 
         .D(\notGate[31]_keep ), .Z(\notGate[32] )) /* synthesis syn_instantiated=1, lut_function=((!D !C !B !A)+(!D !C !B A)+(!D !C B !A)+(!D !C B A)+(!D C !B !A)+(!D C !B A)+(!D C B !A)+(!D C B A)), LSE_LINE_FILE_ID=3, LSE_LCOL=13, LSE_RCOL=44, LSE_LLINE=32, LSE_RLINE=32 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(11[2:53])
    defparam I1.init = 16'b0000000011111111;
    
endmodule
//
// Verilog Description of module inverter_U744
//

module inverter_U744 (\notGate[328]_keep , \notGate[329] ) /* synthesis syn_module_defined=1 */ ;
    input \notGate[328]_keep ;
    output \notGate[329] ;
    
    wire \notGate[328]_keep  /* synthesis alspreserve=1 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(25[15:22])
    
    LUT4 I1 (.A(\notGate[328]_keep ), .B(\notGate[328]_keep ), .C(\notGate[328]_keep ), 
         .D(\notGate[328]_keep ), .Z(\notGate[329] )) /* synthesis syn_instantiated=1, lut_function=((!D !C !B !A)+(!D !C !B A)+(!D !C B !A)+(!D !C B A)+(!D C !B !A)+(!D C !B A)+(!D C B !A)+(!D C B A)), LSE_LINE_FILE_ID=3, LSE_LCOL=13, LSE_RCOL=44, LSE_LLINE=32, LSE_RLINE=32 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(11[2:53])
    defparam I1.init = 16'b0000000011111111;
    
endmodule
//
// Verilog Description of module inverter_U745
//

module inverter_U745 (\notGate[327]_keep , \notGate[328] ) /* synthesis syn_module_defined=1 */ ;
    input \notGate[327]_keep ;
    output \notGate[328] ;
    
    wire \notGate[327]_keep  /* synthesis alspreserve=1 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(25[15:22])
    
    LUT4 I1 (.A(\notGate[327]_keep ), .B(\notGate[327]_keep ), .C(\notGate[327]_keep ), 
         .D(\notGate[327]_keep ), .Z(\notGate[328] )) /* synthesis syn_instantiated=1, lut_function=((!D !C !B !A)+(!D !C !B A)+(!D !C B !A)+(!D !C B A)+(!D C !B !A)+(!D C !B A)+(!D C B !A)+(!D C B A)), LSE_LINE_FILE_ID=3, LSE_LCOL=13, LSE_RCOL=44, LSE_LLINE=32, LSE_RLINE=32 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(11[2:53])
    defparam I1.init = 16'b0000000011111111;
    
endmodule
//
// Verilog Description of module inverter_U746
//

module inverter_U746 (\notGate[326]_keep , \notGate[327] ) /* synthesis syn_module_defined=1 */ ;
    input \notGate[326]_keep ;
    output \notGate[327] ;
    
    wire \notGate[326]_keep  /* synthesis alspreserve=1 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(25[15:22])
    
    LUT4 I1 (.A(\notGate[326]_keep ), .B(\notGate[326]_keep ), .C(\notGate[326]_keep ), 
         .D(\notGate[326]_keep ), .Z(\notGate[327] )) /* synthesis syn_instantiated=1, lut_function=((!D !C !B !A)+(!D !C !B A)+(!D !C B !A)+(!D !C B A)+(!D C !B !A)+(!D C !B A)+(!D C B !A)+(!D C B A)), LSE_LINE_FILE_ID=3, LSE_LCOL=13, LSE_RCOL=44, LSE_LLINE=32, LSE_RLINE=32 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(11[2:53])
    defparam I1.init = 16'b0000000011111111;
    
endmodule
//
// Verilog Description of module inverter_U747
//

module inverter_U747 (\notGate[325]_keep , \notGate[326] ) /* synthesis syn_module_defined=1 */ ;
    input \notGate[325]_keep ;
    output \notGate[326] ;
    
    wire \notGate[325]_keep  /* synthesis alspreserve=1 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(25[15:22])
    
    LUT4 I1 (.A(\notGate[325]_keep ), .B(\notGate[325]_keep ), .C(\notGate[325]_keep ), 
         .D(\notGate[325]_keep ), .Z(\notGate[326] )) /* synthesis syn_instantiated=1, lut_function=((!D !C !B !A)+(!D !C !B A)+(!D !C B !A)+(!D !C B A)+(!D C !B !A)+(!D C !B A)+(!D C B !A)+(!D C B A)), LSE_LINE_FILE_ID=3, LSE_LCOL=13, LSE_RCOL=44, LSE_LLINE=32, LSE_RLINE=32 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(11[2:53])
    defparam I1.init = 16'b0000000011111111;
    
endmodule
//
// Verilog Description of module inverter_U748
//

module inverter_U748 (\notGate[324]_keep , \notGate[325] ) /* synthesis syn_module_defined=1 */ ;
    input \notGate[324]_keep ;
    output \notGate[325] ;
    
    wire \notGate[324]_keep  /* synthesis alspreserve=1 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(25[15:22])
    
    LUT4 I1 (.A(\notGate[324]_keep ), .B(\notGate[324]_keep ), .C(\notGate[324]_keep ), 
         .D(\notGate[324]_keep ), .Z(\notGate[325] )) /* synthesis syn_instantiated=1, lut_function=((!D !C !B !A)+(!D !C !B A)+(!D !C B !A)+(!D !C B A)+(!D C !B !A)+(!D C !B A)+(!D C B !A)+(!D C B A)), LSE_LINE_FILE_ID=3, LSE_LCOL=13, LSE_RCOL=44, LSE_LLINE=32, LSE_RLINE=32 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(11[2:53])
    defparam I1.init = 16'b0000000011111111;
    
endmodule
//
// Verilog Description of module inverter_U749
//

module inverter_U749 (\notGate[323]_keep , \notGate[324] ) /* synthesis syn_module_defined=1 */ ;
    input \notGate[323]_keep ;
    output \notGate[324] ;
    
    wire \notGate[323]_keep  /* synthesis alspreserve=1 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(25[15:22])
    
    LUT4 I1 (.A(\notGate[323]_keep ), .B(\notGate[323]_keep ), .C(\notGate[323]_keep ), 
         .D(\notGate[323]_keep ), .Z(\notGate[324] )) /* synthesis syn_instantiated=1, lut_function=((!D !C !B !A)+(!D !C !B A)+(!D !C B !A)+(!D !C B A)+(!D C !B !A)+(!D C !B A)+(!D C B !A)+(!D C B A)), LSE_LINE_FILE_ID=3, LSE_LCOL=13, LSE_RCOL=44, LSE_LLINE=32, LSE_RLINE=32 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(11[2:53])
    defparam I1.init = 16'b0000000011111111;
    
endmodule
//
// Verilog Description of module inverter_U750
//

module inverter_U750 (\notGate[322]_keep , \notGate[323] ) /* synthesis syn_module_defined=1 */ ;
    input \notGate[322]_keep ;
    output \notGate[323] ;
    
    wire \notGate[322]_keep  /* synthesis alspreserve=1 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(25[15:22])
    
    LUT4 I1 (.A(\notGate[322]_keep ), .B(\notGate[322]_keep ), .C(\notGate[322]_keep ), 
         .D(\notGate[322]_keep ), .Z(\notGate[323] )) /* synthesis syn_instantiated=1, lut_function=((!D !C !B !A)+(!D !C !B A)+(!D !C B !A)+(!D !C B A)+(!D C !B !A)+(!D C !B A)+(!D C B !A)+(!D C B A)), LSE_LINE_FILE_ID=3, LSE_LCOL=13, LSE_RCOL=44, LSE_LLINE=32, LSE_RLINE=32 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(11[2:53])
    defparam I1.init = 16'b0000000011111111;
    
endmodule
//
// Verilog Description of module inverter_U751
//

module inverter_U751 (\notGate[321]_keep , \notGate[322] ) /* synthesis syn_module_defined=1 */ ;
    input \notGate[321]_keep ;
    output \notGate[322] ;
    
    wire \notGate[321]_keep  /* synthesis alspreserve=1 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(25[15:22])
    
    LUT4 I1 (.A(\notGate[321]_keep ), .B(\notGate[321]_keep ), .C(\notGate[321]_keep ), 
         .D(\notGate[321]_keep ), .Z(\notGate[322] )) /* synthesis syn_instantiated=1, lut_function=((!D !C !B !A)+(!D !C !B A)+(!D !C B !A)+(!D !C B A)+(!D C !B !A)+(!D C !B A)+(!D C B !A)+(!D C B A)), LSE_LINE_FILE_ID=3, LSE_LCOL=13, LSE_RCOL=44, LSE_LLINE=32, LSE_RLINE=32 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(11[2:53])
    defparam I1.init = 16'b0000000011111111;
    
endmodule
//
// Verilog Description of module inverter_U752
//

module inverter_U752 (\notGate[320]_keep , \notGate[321] ) /* synthesis syn_module_defined=1 */ ;
    input \notGate[320]_keep ;
    output \notGate[321] ;
    
    wire \notGate[320]_keep  /* synthesis alspreserve=1 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(25[15:22])
    
    LUT4 I1 (.A(\notGate[320]_keep ), .B(\notGate[320]_keep ), .C(\notGate[320]_keep ), 
         .D(\notGate[320]_keep ), .Z(\notGate[321] )) /* synthesis syn_instantiated=1, lut_function=((!D !C !B !A)+(!D !C !B A)+(!D !C B !A)+(!D !C B A)+(!D C !B !A)+(!D C !B A)+(!D C B !A)+(!D C B A)), LSE_LINE_FILE_ID=3, LSE_LCOL=13, LSE_RCOL=44, LSE_LLINE=32, LSE_RLINE=32 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(11[2:53])
    defparam I1.init = 16'b0000000011111111;
    
endmodule
//
// Verilog Description of module inverter_U753
//

module inverter_U753 (\notGate[319]_keep , \notGate[320] ) /* synthesis syn_module_defined=1 */ ;
    input \notGate[319]_keep ;
    output \notGate[320] ;
    
    wire \notGate[319]_keep  /* synthesis alspreserve=1 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(25[15:22])
    
    LUT4 I1 (.A(\notGate[319]_keep ), .B(\notGate[319]_keep ), .C(\notGate[319]_keep ), 
         .D(\notGate[319]_keep ), .Z(\notGate[320] )) /* synthesis syn_instantiated=1, lut_function=((!D !C !B !A)+(!D !C !B A)+(!D !C B !A)+(!D !C B A)+(!D C !B !A)+(!D C !B A)+(!D C B !A)+(!D C B A)), LSE_LINE_FILE_ID=3, LSE_LCOL=13, LSE_RCOL=44, LSE_LLINE=32, LSE_RLINE=32 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(11[2:53])
    defparam I1.init = 16'b0000000011111111;
    
endmodule
//
// Verilog Description of module inverter_U754
//

module inverter_U754 (\notGate[30]_keep , \notGate[31] ) /* synthesis syn_module_defined=1 */ ;
    input \notGate[30]_keep ;
    output \notGate[31] ;
    
    wire \notGate[30]_keep  /* synthesis alspreserve=1 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(25[15:22])
    
    LUT4 I1 (.A(\notGate[30]_keep ), .B(\notGate[30]_keep ), .C(\notGate[30]_keep ), 
         .D(\notGate[30]_keep ), .Z(\notGate[31] )) /* synthesis syn_instantiated=1, lut_function=((!D !C !B !A)+(!D !C !B A)+(!D !C B !A)+(!D !C B A)+(!D C !B !A)+(!D C !B A)+(!D C B !A)+(!D C B A)), LSE_LINE_FILE_ID=3, LSE_LCOL=13, LSE_RCOL=44, LSE_LLINE=32, LSE_RLINE=32 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(11[2:53])
    defparam I1.init = 16'b0000000011111111;
    
endmodule
//
// Verilog Description of module inverter_U755
//

module inverter_U755 (\notGate[318]_keep , \notGate[319] ) /* synthesis syn_module_defined=1 */ ;
    input \notGate[318]_keep ;
    output \notGate[319] ;
    
    wire \notGate[318]_keep  /* synthesis alspreserve=1 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(25[15:22])
    
    LUT4 I1 (.A(\notGate[318]_keep ), .B(\notGate[318]_keep ), .C(\notGate[318]_keep ), 
         .D(\notGate[318]_keep ), .Z(\notGate[319] )) /* synthesis syn_instantiated=1, lut_function=((!D !C !B !A)+(!D !C !B A)+(!D !C B !A)+(!D !C B A)+(!D C !B !A)+(!D C !B A)+(!D C B !A)+(!D C B A)), LSE_LINE_FILE_ID=3, LSE_LCOL=13, LSE_RCOL=44, LSE_LLINE=32, LSE_RLINE=32 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(11[2:53])
    defparam I1.init = 16'b0000000011111111;
    
endmodule
//
// Verilog Description of module inverter_U756
//

module inverter_U756 (\notGate[317]_keep , \notGate[318] ) /* synthesis syn_module_defined=1 */ ;
    input \notGate[317]_keep ;
    output \notGate[318] ;
    
    wire \notGate[317]_keep  /* synthesis alspreserve=1 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(25[15:22])
    
    LUT4 I1 (.A(\notGate[317]_keep ), .B(\notGate[317]_keep ), .C(\notGate[317]_keep ), 
         .D(\notGate[317]_keep ), .Z(\notGate[318] )) /* synthesis syn_instantiated=1, lut_function=((!D !C !B !A)+(!D !C !B A)+(!D !C B !A)+(!D !C B A)+(!D C !B !A)+(!D C !B A)+(!D C B !A)+(!D C B A)), LSE_LINE_FILE_ID=3, LSE_LCOL=13, LSE_RCOL=44, LSE_LLINE=32, LSE_RLINE=32 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(11[2:53])
    defparam I1.init = 16'b0000000011111111;
    
endmodule
//
// Verilog Description of module inverter_U757
//

module inverter_U757 (\notGate[316]_keep , \notGate[317] ) /* synthesis syn_module_defined=1 */ ;
    input \notGate[316]_keep ;
    output \notGate[317] ;
    
    wire \notGate[316]_keep  /* synthesis alspreserve=1 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(25[15:22])
    
    LUT4 I1 (.A(\notGate[316]_keep ), .B(\notGate[316]_keep ), .C(\notGate[316]_keep ), 
         .D(\notGate[316]_keep ), .Z(\notGate[317] )) /* synthesis syn_instantiated=1, lut_function=((!D !C !B !A)+(!D !C !B A)+(!D !C B !A)+(!D !C B A)+(!D C !B !A)+(!D C !B A)+(!D C B !A)+(!D C B A)), LSE_LINE_FILE_ID=3, LSE_LCOL=13, LSE_RCOL=44, LSE_LLINE=32, LSE_RLINE=32 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(11[2:53])
    defparam I1.init = 16'b0000000011111111;
    
endmodule
//
// Verilog Description of module inverter_U758
//

module inverter_U758 (\notGate[315]_keep , \notGate[316] ) /* synthesis syn_module_defined=1 */ ;
    input \notGate[315]_keep ;
    output \notGate[316] ;
    
    wire \notGate[315]_keep  /* synthesis alspreserve=1 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(25[15:22])
    
    LUT4 I1 (.A(\notGate[315]_keep ), .B(\notGate[315]_keep ), .C(\notGate[315]_keep ), 
         .D(\notGate[315]_keep ), .Z(\notGate[316] )) /* synthesis syn_instantiated=1, lut_function=((!D !C !B !A)+(!D !C !B A)+(!D !C B !A)+(!D !C B A)+(!D C !B !A)+(!D C !B A)+(!D C B !A)+(!D C B A)), LSE_LINE_FILE_ID=3, LSE_LCOL=13, LSE_RCOL=44, LSE_LLINE=32, LSE_RLINE=32 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(11[2:53])
    defparam I1.init = 16'b0000000011111111;
    
endmodule
//
// Verilog Description of module inverter_U759
//

module inverter_U759 (\notGate[314]_keep , \notGate[315] ) /* synthesis syn_module_defined=1 */ ;
    input \notGate[314]_keep ;
    output \notGate[315] ;
    
    wire \notGate[314]_keep  /* synthesis alspreserve=1 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(25[15:22])
    
    LUT4 I1 (.A(\notGate[314]_keep ), .B(\notGate[314]_keep ), .C(\notGate[314]_keep ), 
         .D(\notGate[314]_keep ), .Z(\notGate[315] )) /* synthesis syn_instantiated=1, lut_function=((!D !C !B !A)+(!D !C !B A)+(!D !C B !A)+(!D !C B A)+(!D C !B !A)+(!D C !B A)+(!D C B !A)+(!D C B A)), LSE_LINE_FILE_ID=3, LSE_LCOL=13, LSE_RCOL=44, LSE_LLINE=32, LSE_RLINE=32 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(11[2:53])
    defparam I1.init = 16'b0000000011111111;
    
endmodule
//
// Verilog Description of module inverter_U760
//

module inverter_U760 (\notGate[313]_keep , \notGate[314] ) /* synthesis syn_module_defined=1 */ ;
    input \notGate[313]_keep ;
    output \notGate[314] ;
    
    wire \notGate[313]_keep  /* synthesis alspreserve=1 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(25[15:22])
    
    LUT4 I1 (.A(\notGate[313]_keep ), .B(\notGate[313]_keep ), .C(\notGate[313]_keep ), 
         .D(\notGate[313]_keep ), .Z(\notGate[314] )) /* synthesis syn_instantiated=1, lut_function=((!D !C !B !A)+(!D !C !B A)+(!D !C B !A)+(!D !C B A)+(!D C !B !A)+(!D C !B A)+(!D C B !A)+(!D C B A)), LSE_LINE_FILE_ID=3, LSE_LCOL=13, LSE_RCOL=44, LSE_LLINE=32, LSE_RLINE=32 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(11[2:53])
    defparam I1.init = 16'b0000000011111111;
    
endmodule
//
// Verilog Description of module inverter_U761
//

module inverter_U761 (\notGate[312]_keep , \notGate[313] ) /* synthesis syn_module_defined=1 */ ;
    input \notGate[312]_keep ;
    output \notGate[313] ;
    
    wire \notGate[312]_keep  /* synthesis alspreserve=1 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(25[15:22])
    
    LUT4 I1 (.A(\notGate[312]_keep ), .B(\notGate[312]_keep ), .C(\notGate[312]_keep ), 
         .D(\notGate[312]_keep ), .Z(\notGate[313] )) /* synthesis syn_instantiated=1, lut_function=((!D !C !B !A)+(!D !C !B A)+(!D !C B !A)+(!D !C B A)+(!D C !B !A)+(!D C !B A)+(!D C B !A)+(!D C B A)), LSE_LINE_FILE_ID=3, LSE_LCOL=13, LSE_RCOL=44, LSE_LLINE=32, LSE_RLINE=32 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(11[2:53])
    defparam I1.init = 16'b0000000011111111;
    
endmodule
//
// Verilog Description of module inverter_U762
//

module inverter_U762 (\notGate[311]_keep , \notGate[312] ) /* synthesis syn_module_defined=1 */ ;
    input \notGate[311]_keep ;
    output \notGate[312] ;
    
    wire \notGate[311]_keep  /* synthesis alspreserve=1 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(25[15:22])
    
    LUT4 I1 (.A(\notGate[311]_keep ), .B(\notGate[311]_keep ), .C(\notGate[311]_keep ), 
         .D(\notGate[311]_keep ), .Z(\notGate[312] )) /* synthesis syn_instantiated=1, lut_function=((!D !C !B !A)+(!D !C !B A)+(!D !C B !A)+(!D !C B A)+(!D C !B !A)+(!D C !B A)+(!D C B !A)+(!D C B A)), LSE_LINE_FILE_ID=3, LSE_LCOL=13, LSE_RCOL=44, LSE_LLINE=32, LSE_RLINE=32 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(11[2:53])
    defparam I1.init = 16'b0000000011111111;
    
endmodule
//
// Verilog Description of module inverter_U763
//

module inverter_U763 (\notGate[310]_keep , \notGate[311] ) /* synthesis syn_module_defined=1 */ ;
    input \notGate[310]_keep ;
    output \notGate[311] ;
    
    wire \notGate[310]_keep  /* synthesis alspreserve=1 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(25[15:22])
    
    LUT4 I1 (.A(\notGate[310]_keep ), .B(\notGate[310]_keep ), .C(\notGate[310]_keep ), 
         .D(\notGate[310]_keep ), .Z(\notGate[311] )) /* synthesis syn_instantiated=1, lut_function=((!D !C !B !A)+(!D !C !B A)+(!D !C B !A)+(!D !C B A)+(!D C !B !A)+(!D C !B A)+(!D C B !A)+(!D C B A)), LSE_LINE_FILE_ID=3, LSE_LCOL=13, LSE_RCOL=44, LSE_LLINE=32, LSE_RLINE=32 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(11[2:53])
    defparam I1.init = 16'b0000000011111111;
    
endmodule
//
// Verilog Description of module inverter_U764
//

module inverter_U764 (\notGate[309]_keep , \notGate[310] ) /* synthesis syn_module_defined=1 */ ;
    input \notGate[309]_keep ;
    output \notGate[310] ;
    
    wire \notGate[309]_keep  /* synthesis alspreserve=1 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(25[15:22])
    
    LUT4 I1 (.A(\notGate[309]_keep ), .B(\notGate[309]_keep ), .C(\notGate[309]_keep ), 
         .D(\notGate[309]_keep ), .Z(\notGate[310] )) /* synthesis syn_instantiated=1, lut_function=((!D !C !B !A)+(!D !C !B A)+(!D !C B !A)+(!D !C B A)+(!D C !B !A)+(!D C !B A)+(!D C B !A)+(!D C B A)), LSE_LINE_FILE_ID=3, LSE_LCOL=13, LSE_RCOL=44, LSE_LLINE=32, LSE_RLINE=32 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(11[2:53])
    defparam I1.init = 16'b0000000011111111;
    
endmodule
//
// Verilog Description of module inverter_U765
//

module inverter_U765 (\notGate[29]_keep , \notGate[30] ) /* synthesis syn_module_defined=1 */ ;
    input \notGate[29]_keep ;
    output \notGate[30] ;
    
    wire \notGate[29]_keep  /* synthesis alspreserve=1 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(25[15:22])
    
    LUT4 I1 (.A(\notGate[29]_keep ), .B(\notGate[29]_keep ), .C(\notGate[29]_keep ), 
         .D(\notGate[29]_keep ), .Z(\notGate[30] )) /* synthesis syn_instantiated=1, lut_function=((!D !C !B !A)+(!D !C !B A)+(!D !C B !A)+(!D !C B A)+(!D C !B !A)+(!D C !B A)+(!D C B !A)+(!D C B A)), LSE_LINE_FILE_ID=3, LSE_LCOL=13, LSE_RCOL=44, LSE_LLINE=32, LSE_RLINE=32 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(11[2:53])
    defparam I1.init = 16'b0000000011111111;
    
endmodule
//
// Verilog Description of module inverter_U766
//

module inverter_U766 (\notGate[308]_keep , \notGate[309] ) /* synthesis syn_module_defined=1 */ ;
    input \notGate[308]_keep ;
    output \notGate[309] ;
    
    wire \notGate[308]_keep  /* synthesis alspreserve=1 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(25[15:22])
    
    LUT4 I1 (.A(\notGate[308]_keep ), .B(\notGate[308]_keep ), .C(\notGate[308]_keep ), 
         .D(\notGate[308]_keep ), .Z(\notGate[309] )) /* synthesis syn_instantiated=1, lut_function=((!D !C !B !A)+(!D !C !B A)+(!D !C B !A)+(!D !C B A)+(!D C !B !A)+(!D C !B A)+(!D C B !A)+(!D C B A)), LSE_LINE_FILE_ID=3, LSE_LCOL=13, LSE_RCOL=44, LSE_LLINE=32, LSE_RLINE=32 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(11[2:53])
    defparam I1.init = 16'b0000000011111111;
    
endmodule
//
// Verilog Description of module inverter_U767
//

module inverter_U767 (\notGate[307]_keep , \notGate[308] ) /* synthesis syn_module_defined=1 */ ;
    input \notGate[307]_keep ;
    output \notGate[308] ;
    
    wire \notGate[307]_keep  /* synthesis alspreserve=1 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(25[15:22])
    
    LUT4 I1 (.A(\notGate[307]_keep ), .B(\notGate[307]_keep ), .C(\notGate[307]_keep ), 
         .D(\notGate[307]_keep ), .Z(\notGate[308] )) /* synthesis syn_instantiated=1, lut_function=((!D !C !B !A)+(!D !C !B A)+(!D !C B !A)+(!D !C B A)+(!D C !B !A)+(!D C !B A)+(!D C B !A)+(!D C B A)), LSE_LINE_FILE_ID=3, LSE_LCOL=13, LSE_RCOL=44, LSE_LLINE=32, LSE_RLINE=32 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(11[2:53])
    defparam I1.init = 16'b0000000011111111;
    
endmodule
//
// Verilog Description of module inverter_U768
//

module inverter_U768 (\notGate[306]_keep , \notGate[307] ) /* synthesis syn_module_defined=1 */ ;
    input \notGate[306]_keep ;
    output \notGate[307] ;
    
    wire \notGate[306]_keep  /* synthesis alspreserve=1 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(25[15:22])
    
    LUT4 I1 (.A(\notGate[306]_keep ), .B(\notGate[306]_keep ), .C(\notGate[306]_keep ), 
         .D(\notGate[306]_keep ), .Z(\notGate[307] )) /* synthesis syn_instantiated=1, lut_function=((!D !C !B !A)+(!D !C !B A)+(!D !C B !A)+(!D !C B A)+(!D C !B !A)+(!D C !B A)+(!D C B !A)+(!D C B A)), LSE_LINE_FILE_ID=3, LSE_LCOL=13, LSE_RCOL=44, LSE_LLINE=32, LSE_RLINE=32 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(11[2:53])
    defparam I1.init = 16'b0000000011111111;
    
endmodule
//
// Verilog Description of module inverter_U769
//

module inverter_U769 (\notGate[305]_keep , \notGate[306] ) /* synthesis syn_module_defined=1 */ ;
    input \notGate[305]_keep ;
    output \notGate[306] ;
    
    wire \notGate[305]_keep  /* synthesis alspreserve=1 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(25[15:22])
    
    LUT4 I1 (.A(\notGate[305]_keep ), .B(\notGate[305]_keep ), .C(\notGate[305]_keep ), 
         .D(\notGate[305]_keep ), .Z(\notGate[306] )) /* synthesis syn_instantiated=1, lut_function=((!D !C !B !A)+(!D !C !B A)+(!D !C B !A)+(!D !C B A)+(!D C !B !A)+(!D C !B A)+(!D C B !A)+(!D C B A)), LSE_LINE_FILE_ID=3, LSE_LCOL=13, LSE_RCOL=44, LSE_LLINE=32, LSE_RLINE=32 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(11[2:53])
    defparam I1.init = 16'b0000000011111111;
    
endmodule
//
// Verilog Description of module inverter_U770
//

module inverter_U770 (\notGate[304]_keep , \notGate[305] ) /* synthesis syn_module_defined=1 */ ;
    input \notGate[304]_keep ;
    output \notGate[305] ;
    
    wire \notGate[304]_keep  /* synthesis alspreserve=1 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(25[15:22])
    
    LUT4 I1 (.A(\notGate[304]_keep ), .B(\notGate[304]_keep ), .C(\notGate[304]_keep ), 
         .D(\notGate[304]_keep ), .Z(\notGate[305] )) /* synthesis syn_instantiated=1, lut_function=((!D !C !B !A)+(!D !C !B A)+(!D !C B !A)+(!D !C B A)+(!D C !B !A)+(!D C !B A)+(!D C B !A)+(!D C B A)), LSE_LINE_FILE_ID=3, LSE_LCOL=13, LSE_RCOL=44, LSE_LLINE=32, LSE_RLINE=32 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(11[2:53])
    defparam I1.init = 16'b0000000011111111;
    
endmodule
//
// Verilog Description of module inverter_U771
//

module inverter_U771 (\notGate[303]_keep , \notGate[304] ) /* synthesis syn_module_defined=1 */ ;
    input \notGate[303]_keep ;
    output \notGate[304] ;
    
    wire \notGate[303]_keep  /* synthesis alspreserve=1 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(25[15:22])
    
    LUT4 I1 (.A(\notGate[303]_keep ), .B(\notGate[303]_keep ), .C(\notGate[303]_keep ), 
         .D(\notGate[303]_keep ), .Z(\notGate[304] )) /* synthesis syn_instantiated=1, lut_function=((!D !C !B !A)+(!D !C !B A)+(!D !C B !A)+(!D !C B A)+(!D C !B !A)+(!D C !B A)+(!D C B !A)+(!D C B A)), LSE_LINE_FILE_ID=3, LSE_LCOL=13, LSE_RCOL=44, LSE_LLINE=32, LSE_RLINE=32 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(11[2:53])
    defparam I1.init = 16'b0000000011111111;
    
endmodule
//
// Verilog Description of module inverter_U772
//

module inverter_U772 (\notGate[302]_keep , \notGate[303] ) /* synthesis syn_module_defined=1 */ ;
    input \notGate[302]_keep ;
    output \notGate[303] ;
    
    wire \notGate[302]_keep  /* synthesis alspreserve=1 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(25[15:22])
    
    LUT4 I1 (.A(\notGate[302]_keep ), .B(\notGate[302]_keep ), .C(\notGate[302]_keep ), 
         .D(\notGate[302]_keep ), .Z(\notGate[303] )) /* synthesis syn_instantiated=1, lut_function=((!D !C !B !A)+(!D !C !B A)+(!D !C B !A)+(!D !C B A)+(!D C !B !A)+(!D C !B A)+(!D C B !A)+(!D C B A)), LSE_LINE_FILE_ID=3, LSE_LCOL=13, LSE_RCOL=44, LSE_LLINE=32, LSE_RLINE=32 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(11[2:53])
    defparam I1.init = 16'b0000000011111111;
    
endmodule
//
// Verilog Description of module inverter_U773
//

module inverter_U773 (\notGate[301]_keep , \notGate[302] ) /* synthesis syn_module_defined=1 */ ;
    input \notGate[301]_keep ;
    output \notGate[302] ;
    
    wire \notGate[301]_keep  /* synthesis alspreserve=1 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(25[15:22])
    
    LUT4 I1 (.A(\notGate[301]_keep ), .B(\notGate[301]_keep ), .C(\notGate[301]_keep ), 
         .D(\notGate[301]_keep ), .Z(\notGate[302] )) /* synthesis syn_instantiated=1, lut_function=((!D !C !B !A)+(!D !C !B A)+(!D !C B !A)+(!D !C B A)+(!D C !B !A)+(!D C !B A)+(!D C B !A)+(!D C B A)), LSE_LINE_FILE_ID=3, LSE_LCOL=13, LSE_RCOL=44, LSE_LLINE=32, LSE_RLINE=32 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(11[2:53])
    defparam I1.init = 16'b0000000011111111;
    
endmodule
//
// Verilog Description of module inverter_U774
//

module inverter_U774 (\notGate[300]_keep , \notGate[301] ) /* synthesis syn_module_defined=1 */ ;
    input \notGate[300]_keep ;
    output \notGate[301] ;
    
    wire \notGate[300]_keep  /* synthesis alspreserve=1 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(25[15:22])
    
    LUT4 I1 (.A(\notGate[300]_keep ), .B(\notGate[300]_keep ), .C(\notGate[300]_keep ), 
         .D(\notGate[300]_keep ), .Z(\notGate[301] )) /* synthesis syn_instantiated=1, lut_function=((!D !C !B !A)+(!D !C !B A)+(!D !C B !A)+(!D !C B A)+(!D C !B !A)+(!D C !B A)+(!D C B !A)+(!D C B A)), LSE_LINE_FILE_ID=3, LSE_LCOL=13, LSE_RCOL=44, LSE_LLINE=32, LSE_RLINE=32 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(11[2:53])
    defparam I1.init = 16'b0000000011111111;
    
endmodule
//
// Verilog Description of module inverter_U775
//

module inverter_U775 (\notGate[299]_keep , \notGate[300] ) /* synthesis syn_module_defined=1 */ ;
    input \notGate[299]_keep ;
    output \notGate[300] ;
    
    wire \notGate[299]_keep  /* synthesis alspreserve=1 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(25[15:22])
    
    LUT4 I1 (.A(\notGate[299]_keep ), .B(\notGate[299]_keep ), .C(\notGate[299]_keep ), 
         .D(\notGate[299]_keep ), .Z(\notGate[300] )) /* synthesis syn_instantiated=1, lut_function=((!D !C !B !A)+(!D !C !B A)+(!D !C B !A)+(!D !C B A)+(!D C !B !A)+(!D C !B A)+(!D C B !A)+(!D C B A)), LSE_LINE_FILE_ID=3, LSE_LCOL=13, LSE_RCOL=44, LSE_LLINE=32, LSE_RLINE=32 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(11[2:53])
    defparam I1.init = 16'b0000000011111111;
    
endmodule
//
// Verilog Description of module inverter_U776
//

module inverter_U776 (\notGate[1]_keep , \notGate[2] ) /* synthesis syn_module_defined=1 */ ;
    input \notGate[1]_keep ;
    output \notGate[2] ;
    
    wire \notGate[1]_keep  /* synthesis alspreserve=1 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(25[15:22])
    
    LUT4 I1 (.A(\notGate[1]_keep ), .B(\notGate[1]_keep ), .C(\notGate[1]_keep ), 
         .D(\notGate[1]_keep ), .Z(\notGate[2] )) /* synthesis syn_instantiated=1, lut_function=((!D !C !B !A)+(!D !C !B A)+(!D !C B !A)+(!D !C B A)+(!D C !B !A)+(!D C !B A)+(!D C B !A)+(!D C B A)), LSE_LINE_FILE_ID=3, LSE_LCOL=13, LSE_RCOL=44, LSE_LLINE=32, LSE_RLINE=32 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(11[2:53])
    defparam I1.init = 16'b0000000011111111;
    
endmodule
//
// Verilog Description of module inverter_U777
//

module inverter_U777 (\notGate[28]_keep , \notGate[29] ) /* synthesis syn_module_defined=1 */ ;
    input \notGate[28]_keep ;
    output \notGate[29] ;
    
    wire \notGate[28]_keep  /* synthesis alspreserve=1 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(25[15:22])
    
    LUT4 I1 (.A(\notGate[28]_keep ), .B(\notGate[28]_keep ), .C(\notGate[28]_keep ), 
         .D(\notGate[28]_keep ), .Z(\notGate[29] )) /* synthesis syn_instantiated=1, lut_function=((!D !C !B !A)+(!D !C !B A)+(!D !C B !A)+(!D !C B A)+(!D C !B !A)+(!D C !B A)+(!D C B !A)+(!D C B A)), LSE_LINE_FILE_ID=3, LSE_LCOL=13, LSE_RCOL=44, LSE_LLINE=32, LSE_RLINE=32 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(11[2:53])
    defparam I1.init = 16'b0000000011111111;
    
endmodule
//
// Verilog Description of module inverter_U778
//

module inverter_U778 (\notGate[298]_keep , \notGate[299] ) /* synthesis syn_module_defined=1 */ ;
    input \notGate[298]_keep ;
    output \notGate[299] ;
    
    wire \notGate[298]_keep  /* synthesis alspreserve=1 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(25[15:22])
    
    LUT4 I1 (.A(\notGate[298]_keep ), .B(\notGate[298]_keep ), .C(\notGate[298]_keep ), 
         .D(\notGate[298]_keep ), .Z(\notGate[299] )) /* synthesis syn_instantiated=1, lut_function=((!D !C !B !A)+(!D !C !B A)+(!D !C B !A)+(!D !C B A)+(!D C !B !A)+(!D C !B A)+(!D C B !A)+(!D C B A)), LSE_LINE_FILE_ID=3, LSE_LCOL=13, LSE_RCOL=44, LSE_LLINE=32, LSE_RLINE=32 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(11[2:53])
    defparam I1.init = 16'b0000000011111111;
    
endmodule
//
// Verilog Description of module inverter_U779
//

module inverter_U779 (\notGate[297]_keep , \notGate[298] ) /* synthesis syn_module_defined=1 */ ;
    input \notGate[297]_keep ;
    output \notGate[298] ;
    
    wire \notGate[297]_keep  /* synthesis alspreserve=1 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(25[15:22])
    
    LUT4 I1 (.A(\notGate[297]_keep ), .B(\notGate[297]_keep ), .C(\notGate[297]_keep ), 
         .D(\notGate[297]_keep ), .Z(\notGate[298] )) /* synthesis syn_instantiated=1, lut_function=((!D !C !B !A)+(!D !C !B A)+(!D !C B !A)+(!D !C B A)+(!D C !B !A)+(!D C !B A)+(!D C B !A)+(!D C B A)), LSE_LINE_FILE_ID=3, LSE_LCOL=13, LSE_RCOL=44, LSE_LLINE=32, LSE_RLINE=32 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(11[2:53])
    defparam I1.init = 16'b0000000011111111;
    
endmodule
//
// Verilog Description of module inverter_U780
//

module inverter_U780 (\notGate[296]_keep , \notGate[297] ) /* synthesis syn_module_defined=1 */ ;
    input \notGate[296]_keep ;
    output \notGate[297] ;
    
    wire \notGate[296]_keep  /* synthesis alspreserve=1 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(25[15:22])
    
    LUT4 I1 (.A(\notGate[296]_keep ), .B(\notGate[296]_keep ), .C(\notGate[296]_keep ), 
         .D(\notGate[296]_keep ), .Z(\notGate[297] )) /* synthesis syn_instantiated=1, lut_function=((!D !C !B !A)+(!D !C !B A)+(!D !C B !A)+(!D !C B A)+(!D C !B !A)+(!D C !B A)+(!D C B !A)+(!D C B A)), LSE_LINE_FILE_ID=3, LSE_LCOL=13, LSE_RCOL=44, LSE_LLINE=32, LSE_RLINE=32 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(11[2:53])
    defparam I1.init = 16'b0000000011111111;
    
endmodule
//
// Verilog Description of module inverter_U781
//

module inverter_U781 (\notGate[295]_keep , \notGate[296] ) /* synthesis syn_module_defined=1 */ ;
    input \notGate[295]_keep ;
    output \notGate[296] ;
    
    wire \notGate[295]_keep  /* synthesis alspreserve=1 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(25[15:22])
    
    LUT4 I1 (.A(\notGate[295]_keep ), .B(\notGate[295]_keep ), .C(\notGate[295]_keep ), 
         .D(\notGate[295]_keep ), .Z(\notGate[296] )) /* synthesis syn_instantiated=1, lut_function=((!D !C !B !A)+(!D !C !B A)+(!D !C B !A)+(!D !C B A)+(!D C !B !A)+(!D C !B A)+(!D C B !A)+(!D C B A)), LSE_LINE_FILE_ID=3, LSE_LCOL=13, LSE_RCOL=44, LSE_LLINE=32, LSE_RLINE=32 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(11[2:53])
    defparam I1.init = 16'b0000000011111111;
    
endmodule
//
// Verilog Description of module inverter_U782
//

module inverter_U782 (\notGate[294]_keep , \notGate[295] ) /* synthesis syn_module_defined=1 */ ;
    input \notGate[294]_keep ;
    output \notGate[295] ;
    
    wire \notGate[294]_keep  /* synthesis alspreserve=1 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(25[15:22])
    
    LUT4 I1 (.A(\notGate[294]_keep ), .B(\notGate[294]_keep ), .C(\notGate[294]_keep ), 
         .D(\notGate[294]_keep ), .Z(\notGate[295] )) /* synthesis syn_instantiated=1, lut_function=((!D !C !B !A)+(!D !C !B A)+(!D !C B !A)+(!D !C B A)+(!D C !B !A)+(!D C !B A)+(!D C B !A)+(!D C B A)), LSE_LINE_FILE_ID=3, LSE_LCOL=13, LSE_RCOL=44, LSE_LLINE=32, LSE_RLINE=32 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(11[2:53])
    defparam I1.init = 16'b0000000011111111;
    
endmodule
//
// Verilog Description of module inverter_U783
//

module inverter_U783 (\notGate[293]_keep , \notGate[294] ) /* synthesis syn_module_defined=1 */ ;
    input \notGate[293]_keep ;
    output \notGate[294] ;
    
    wire \notGate[293]_keep  /* synthesis alspreserve=1 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(25[15:22])
    
    LUT4 I1 (.A(\notGate[293]_keep ), .B(\notGate[293]_keep ), .C(\notGate[293]_keep ), 
         .D(\notGate[293]_keep ), .Z(\notGate[294] )) /* synthesis syn_instantiated=1, lut_function=((!D !C !B !A)+(!D !C !B A)+(!D !C B !A)+(!D !C B A)+(!D C !B !A)+(!D C !B A)+(!D C B !A)+(!D C B A)), LSE_LINE_FILE_ID=3, LSE_LCOL=13, LSE_RCOL=44, LSE_LLINE=32, LSE_RLINE=32 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(11[2:53])
    defparam I1.init = 16'b0000000011111111;
    
endmodule
//
// Verilog Description of module inverter_U784
//

module inverter_U784 (\notGate[292]_keep , \notGate[293] ) /* synthesis syn_module_defined=1 */ ;
    input \notGate[292]_keep ;
    output \notGate[293] ;
    
    wire \notGate[292]_keep  /* synthesis alspreserve=1 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(25[15:22])
    
    LUT4 I1 (.A(\notGate[292]_keep ), .B(\notGate[292]_keep ), .C(\notGate[292]_keep ), 
         .D(\notGate[292]_keep ), .Z(\notGate[293] )) /* synthesis syn_instantiated=1, lut_function=((!D !C !B !A)+(!D !C !B A)+(!D !C B !A)+(!D !C B A)+(!D C !B !A)+(!D C !B A)+(!D C B !A)+(!D C B A)), LSE_LINE_FILE_ID=3, LSE_LCOL=13, LSE_RCOL=44, LSE_LLINE=32, LSE_RLINE=32 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(11[2:53])
    defparam I1.init = 16'b0000000011111111;
    
endmodule
//
// Verilog Description of module inverter_U785
//

module inverter_U785 (\notGate[291]_keep , \notGate[292] ) /* synthesis syn_module_defined=1 */ ;
    input \notGate[291]_keep ;
    output \notGate[292] ;
    
    wire \notGate[291]_keep  /* synthesis alspreserve=1 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(25[15:22])
    
    LUT4 I1 (.A(\notGate[291]_keep ), .B(\notGate[291]_keep ), .C(\notGate[291]_keep ), 
         .D(\notGate[291]_keep ), .Z(\notGate[292] )) /* synthesis syn_instantiated=1, lut_function=((!D !C !B !A)+(!D !C !B A)+(!D !C B !A)+(!D !C B A)+(!D C !B !A)+(!D C !B A)+(!D C B !A)+(!D C B A)), LSE_LINE_FILE_ID=3, LSE_LCOL=13, LSE_RCOL=44, LSE_LLINE=32, LSE_RLINE=32 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(11[2:53])
    defparam I1.init = 16'b0000000011111111;
    
endmodule
//
// Verilog Description of module inverter_U786
//

module inverter_U786 (\notGate[290]_keep , \notGate[291] ) /* synthesis syn_module_defined=1 */ ;
    input \notGate[290]_keep ;
    output \notGate[291] ;
    
    wire \notGate[290]_keep  /* synthesis alspreserve=1 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(25[15:22])
    
    LUT4 I1 (.A(\notGate[290]_keep ), .B(\notGate[290]_keep ), .C(\notGate[290]_keep ), 
         .D(\notGate[290]_keep ), .Z(\notGate[291] )) /* synthesis syn_instantiated=1, lut_function=((!D !C !B !A)+(!D !C !B A)+(!D !C B !A)+(!D !C B A)+(!D C !B !A)+(!D C !B A)+(!D C B !A)+(!D C B A)), LSE_LINE_FILE_ID=3, LSE_LCOL=13, LSE_RCOL=44, LSE_LLINE=32, LSE_RLINE=32 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(11[2:53])
    defparam I1.init = 16'b0000000011111111;
    
endmodule
//
// Verilog Description of module inverter_U787
//

module inverter_U787 (\notGate[289]_keep , \notGate[290] ) /* synthesis syn_module_defined=1 */ ;
    input \notGate[289]_keep ;
    output \notGate[290] ;
    
    wire \notGate[289]_keep  /* synthesis alspreserve=1 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(25[15:22])
    
    LUT4 I1 (.A(\notGate[289]_keep ), .B(\notGate[289]_keep ), .C(\notGate[289]_keep ), 
         .D(\notGate[289]_keep ), .Z(\notGate[290] )) /* synthesis syn_instantiated=1, lut_function=((!D !C !B !A)+(!D !C !B A)+(!D !C B !A)+(!D !C B A)+(!D C !B !A)+(!D C !B A)+(!D C B !A)+(!D C B A)), LSE_LINE_FILE_ID=3, LSE_LCOL=13, LSE_RCOL=44, LSE_LLINE=32, LSE_RLINE=32 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(11[2:53])
    defparam I1.init = 16'b0000000011111111;
    
endmodule
//
// Verilog Description of module inverter_U788
//

module inverter_U788 (\notGate[27]_keep , \notGate[28] ) /* synthesis syn_module_defined=1 */ ;
    input \notGate[27]_keep ;
    output \notGate[28] ;
    
    wire \notGate[27]_keep  /* synthesis alspreserve=1 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(25[15:22])
    
    LUT4 I1 (.A(\notGate[27]_keep ), .B(\notGate[27]_keep ), .C(\notGate[27]_keep ), 
         .D(\notGate[27]_keep ), .Z(\notGate[28] )) /* synthesis syn_instantiated=1, lut_function=((!D !C !B !A)+(!D !C !B A)+(!D !C B !A)+(!D !C B A)+(!D C !B !A)+(!D C !B A)+(!D C B !A)+(!D C B A)), LSE_LINE_FILE_ID=3, LSE_LCOL=13, LSE_RCOL=44, LSE_LLINE=32, LSE_RLINE=32 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(11[2:53])
    defparam I1.init = 16'b0000000011111111;
    
endmodule
//
// Verilog Description of module inverter_U789
//

module inverter_U789 (\notGate[288]_keep , \notGate[289] ) /* synthesis syn_module_defined=1 */ ;
    input \notGate[288]_keep ;
    output \notGate[289] ;
    
    wire \notGate[288]_keep  /* synthesis alspreserve=1 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(25[15:22])
    
    LUT4 I1 (.A(\notGate[288]_keep ), .B(\notGate[288]_keep ), .C(\notGate[288]_keep ), 
         .D(\notGate[288]_keep ), .Z(\notGate[289] )) /* synthesis syn_instantiated=1, lut_function=((!D !C !B !A)+(!D !C !B A)+(!D !C B !A)+(!D !C B A)+(!D C !B !A)+(!D C !B A)+(!D C B !A)+(!D C B A)), LSE_LINE_FILE_ID=3, LSE_LCOL=13, LSE_RCOL=44, LSE_LLINE=32, LSE_RLINE=32 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(11[2:53])
    defparam I1.init = 16'b0000000011111111;
    
endmodule
//
// Verilog Description of module inverter_U790
//

module inverter_U790 (\notGate[287]_keep , \notGate[288] ) /* synthesis syn_module_defined=1 */ ;
    input \notGate[287]_keep ;
    output \notGate[288] ;
    
    wire \notGate[287]_keep  /* synthesis alspreserve=1 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(25[15:22])
    
    LUT4 I1 (.A(\notGate[287]_keep ), .B(\notGate[287]_keep ), .C(\notGate[287]_keep ), 
         .D(\notGate[287]_keep ), .Z(\notGate[288] )) /* synthesis syn_instantiated=1, lut_function=((!D !C !B !A)+(!D !C !B A)+(!D !C B !A)+(!D !C B A)+(!D C !B !A)+(!D C !B A)+(!D C B !A)+(!D C B A)), LSE_LINE_FILE_ID=3, LSE_LCOL=13, LSE_RCOL=44, LSE_LLINE=32, LSE_RLINE=32 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(11[2:53])
    defparam I1.init = 16'b0000000011111111;
    
endmodule
//
// Verilog Description of module inverter_U791
//

module inverter_U791 (\notGate[286]_keep , \notGate[287] ) /* synthesis syn_module_defined=1 */ ;
    input \notGate[286]_keep ;
    output \notGate[287] ;
    
    wire \notGate[286]_keep  /* synthesis alspreserve=1 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(25[15:22])
    
    LUT4 I1 (.A(\notGate[286]_keep ), .B(\notGate[286]_keep ), .C(\notGate[286]_keep ), 
         .D(\notGate[286]_keep ), .Z(\notGate[287] )) /* synthesis syn_instantiated=1, lut_function=((!D !C !B !A)+(!D !C !B A)+(!D !C B !A)+(!D !C B A)+(!D C !B !A)+(!D C !B A)+(!D C B !A)+(!D C B A)), LSE_LINE_FILE_ID=3, LSE_LCOL=13, LSE_RCOL=44, LSE_LLINE=32, LSE_RLINE=32 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(11[2:53])
    defparam I1.init = 16'b0000000011111111;
    
endmodule
//
// Verilog Description of module inverter_U792
//

module inverter_U792 (\notGate[285]_keep , \notGate[286] ) /* synthesis syn_module_defined=1 */ ;
    input \notGate[285]_keep ;
    output \notGate[286] ;
    
    wire \notGate[285]_keep  /* synthesis alspreserve=1 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(25[15:22])
    
    LUT4 I1 (.A(\notGate[285]_keep ), .B(\notGate[285]_keep ), .C(\notGate[285]_keep ), 
         .D(\notGate[285]_keep ), .Z(\notGate[286] )) /* synthesis syn_instantiated=1, lut_function=((!D !C !B !A)+(!D !C !B A)+(!D !C B !A)+(!D !C B A)+(!D C !B !A)+(!D C !B A)+(!D C B !A)+(!D C B A)), LSE_LINE_FILE_ID=3, LSE_LCOL=13, LSE_RCOL=44, LSE_LLINE=32, LSE_RLINE=32 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(11[2:53])
    defparam I1.init = 16'b0000000011111111;
    
endmodule
//
// Verilog Description of module inverter_U793
//

module inverter_U793 (\notGate[284]_keep , \notGate[285] ) /* synthesis syn_module_defined=1 */ ;
    input \notGate[284]_keep ;
    output \notGate[285] ;
    
    wire \notGate[284]_keep  /* synthesis alspreserve=1 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(25[15:22])
    
    LUT4 I1 (.A(\notGate[284]_keep ), .B(\notGate[284]_keep ), .C(\notGate[284]_keep ), 
         .D(\notGate[284]_keep ), .Z(\notGate[285] )) /* synthesis syn_instantiated=1, lut_function=((!D !C !B !A)+(!D !C !B A)+(!D !C B !A)+(!D !C B A)+(!D C !B !A)+(!D C !B A)+(!D C B !A)+(!D C B A)), LSE_LINE_FILE_ID=3, LSE_LCOL=13, LSE_RCOL=44, LSE_LLINE=32, LSE_RLINE=32 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(11[2:53])
    defparam I1.init = 16'b0000000011111111;
    
endmodule
//
// Verilog Description of module inverter_U794
//

module inverter_U794 (\notGate[283]_keep , \notGate[284] ) /* synthesis syn_module_defined=1 */ ;
    input \notGate[283]_keep ;
    output \notGate[284] ;
    
    wire \notGate[283]_keep  /* synthesis alspreserve=1 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(25[15:22])
    
    LUT4 I1 (.A(\notGate[283]_keep ), .B(\notGate[283]_keep ), .C(\notGate[283]_keep ), 
         .D(\notGate[283]_keep ), .Z(\notGate[284] )) /* synthesis syn_instantiated=1, lut_function=((!D !C !B !A)+(!D !C !B A)+(!D !C B !A)+(!D !C B A)+(!D C !B !A)+(!D C !B A)+(!D C B !A)+(!D C B A)), LSE_LINE_FILE_ID=3, LSE_LCOL=13, LSE_RCOL=44, LSE_LLINE=32, LSE_RLINE=32 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(11[2:53])
    defparam I1.init = 16'b0000000011111111;
    
endmodule
//
// Verilog Description of module inverter_U795
//

module inverter_U795 (\notGate[282]_keep , \notGate[283] ) /* synthesis syn_module_defined=1 */ ;
    input \notGate[282]_keep ;
    output \notGate[283] ;
    
    wire \notGate[282]_keep  /* synthesis alspreserve=1 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(25[15:22])
    
    LUT4 I1 (.A(\notGate[282]_keep ), .B(\notGate[282]_keep ), .C(\notGate[282]_keep ), 
         .D(\notGate[282]_keep ), .Z(\notGate[283] )) /* synthesis syn_instantiated=1, lut_function=((!D !C !B !A)+(!D !C !B A)+(!D !C B !A)+(!D !C B A)+(!D C !B !A)+(!D C !B A)+(!D C B !A)+(!D C B A)), LSE_LINE_FILE_ID=3, LSE_LCOL=13, LSE_RCOL=44, LSE_LLINE=32, LSE_RLINE=32 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(11[2:53])
    defparam I1.init = 16'b0000000011111111;
    
endmodule
//
// Verilog Description of module inverter_U796
//

module inverter_U796 (\notGate[281]_keep , \notGate[282] ) /* synthesis syn_module_defined=1 */ ;
    input \notGate[281]_keep ;
    output \notGate[282] ;
    
    wire \notGate[281]_keep  /* synthesis alspreserve=1 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(25[15:22])
    
    LUT4 I1 (.A(\notGate[281]_keep ), .B(\notGate[281]_keep ), .C(\notGate[281]_keep ), 
         .D(\notGate[281]_keep ), .Z(\notGate[282] )) /* synthesis syn_instantiated=1, lut_function=((!D !C !B !A)+(!D !C !B A)+(!D !C B !A)+(!D !C B A)+(!D C !B !A)+(!D C !B A)+(!D C B !A)+(!D C B A)), LSE_LINE_FILE_ID=3, LSE_LCOL=13, LSE_RCOL=44, LSE_LLINE=32, LSE_RLINE=32 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(11[2:53])
    defparam I1.init = 16'b0000000011111111;
    
endmodule
//
// Verilog Description of module inverter_U797
//

module inverter_U797 (\notGate[280]_keep , \notGate[281] ) /* synthesis syn_module_defined=1 */ ;
    input \notGate[280]_keep ;
    output \notGate[281] ;
    
    wire \notGate[280]_keep  /* synthesis alspreserve=1 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(25[15:22])
    
    LUT4 I1 (.A(\notGate[280]_keep ), .B(\notGate[280]_keep ), .C(\notGate[280]_keep ), 
         .D(\notGate[280]_keep ), .Z(\notGate[281] )) /* synthesis syn_instantiated=1, lut_function=((!D !C !B !A)+(!D !C !B A)+(!D !C B !A)+(!D !C B A)+(!D C !B !A)+(!D C !B A)+(!D C B !A)+(!D C B A)), LSE_LINE_FILE_ID=3, LSE_LCOL=13, LSE_RCOL=44, LSE_LLINE=32, LSE_RLINE=32 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(11[2:53])
    defparam I1.init = 16'b0000000011111111;
    
endmodule
//
// Verilog Description of module inverter_U798
//

module inverter_U798 (\notGate[279]_keep , \notGate[280] ) /* synthesis syn_module_defined=1 */ ;
    input \notGate[279]_keep ;
    output \notGate[280] ;
    
    wire \notGate[279]_keep  /* synthesis alspreserve=1 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(25[15:22])
    
    LUT4 I1 (.A(\notGate[279]_keep ), .B(\notGate[279]_keep ), .C(\notGate[279]_keep ), 
         .D(\notGate[279]_keep ), .Z(\notGate[280] )) /* synthesis syn_instantiated=1, lut_function=((!D !C !B !A)+(!D !C !B A)+(!D !C B !A)+(!D !C B A)+(!D C !B !A)+(!D C !B A)+(!D C B !A)+(!D C B A)), LSE_LINE_FILE_ID=3, LSE_LCOL=13, LSE_RCOL=44, LSE_LLINE=32, LSE_RLINE=32 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(11[2:53])
    defparam I1.init = 16'b0000000011111111;
    
endmodule
//
// Verilog Description of module inverter_U799
//

module inverter_U799 (\notGate[26]_keep , \notGate[27] ) /* synthesis syn_module_defined=1 */ ;
    input \notGate[26]_keep ;
    output \notGate[27] ;
    
    wire \notGate[26]_keep  /* synthesis alspreserve=1 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(25[15:22])
    
    LUT4 I1 (.A(\notGate[26]_keep ), .B(\notGate[26]_keep ), .C(\notGate[26]_keep ), 
         .D(\notGate[26]_keep ), .Z(\notGate[27] )) /* synthesis syn_instantiated=1, lut_function=((!D !C !B !A)+(!D !C !B A)+(!D !C B !A)+(!D !C B A)+(!D C !B !A)+(!D C !B A)+(!D C B !A)+(!D C B A)), LSE_LINE_FILE_ID=3, LSE_LCOL=13, LSE_RCOL=44, LSE_LLINE=32, LSE_RLINE=32 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(11[2:53])
    defparam I1.init = 16'b0000000011111111;
    
endmodule
//
// Verilog Description of module inverter_U800
//

module inverter_U800 (\notGate[278]_keep , \notGate[279] ) /* synthesis syn_module_defined=1 */ ;
    input \notGate[278]_keep ;
    output \notGate[279] ;
    
    wire \notGate[278]_keep  /* synthesis alspreserve=1 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(25[15:22])
    
    LUT4 I1 (.A(\notGate[278]_keep ), .B(\notGate[278]_keep ), .C(\notGate[278]_keep ), 
         .D(\notGate[278]_keep ), .Z(\notGate[279] )) /* synthesis syn_instantiated=1, lut_function=((!D !C !B !A)+(!D !C !B A)+(!D !C B !A)+(!D !C B A)+(!D C !B !A)+(!D C !B A)+(!D C B !A)+(!D C B A)), LSE_LINE_FILE_ID=3, LSE_LCOL=13, LSE_RCOL=44, LSE_LLINE=32, LSE_RLINE=32 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(11[2:53])
    defparam I1.init = 16'b0000000011111111;
    
endmodule
//
// Verilog Description of module inverter_U801
//

module inverter_U801 (\notGate[277]_keep , \notGate[278] ) /* synthesis syn_module_defined=1 */ ;
    input \notGate[277]_keep ;
    output \notGate[278] ;
    
    wire \notGate[277]_keep  /* synthesis alspreserve=1 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(25[15:22])
    
    LUT4 I1 (.A(\notGate[277]_keep ), .B(\notGate[277]_keep ), .C(\notGate[277]_keep ), 
         .D(\notGate[277]_keep ), .Z(\notGate[278] )) /* synthesis syn_instantiated=1, lut_function=((!D !C !B !A)+(!D !C !B A)+(!D !C B !A)+(!D !C B A)+(!D C !B !A)+(!D C !B A)+(!D C B !A)+(!D C B A)), LSE_LINE_FILE_ID=3, LSE_LCOL=13, LSE_RCOL=44, LSE_LLINE=32, LSE_RLINE=32 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(11[2:53])
    defparam I1.init = 16'b0000000011111111;
    
endmodule
//
// Verilog Description of module inverter_U802
//

module inverter_U802 (\notGate[276]_keep , \notGate[277] ) /* synthesis syn_module_defined=1 */ ;
    input \notGate[276]_keep ;
    output \notGate[277] ;
    
    wire \notGate[276]_keep  /* synthesis alspreserve=1 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(25[15:22])
    
    LUT4 I1 (.A(\notGate[276]_keep ), .B(\notGate[276]_keep ), .C(\notGate[276]_keep ), 
         .D(\notGate[276]_keep ), .Z(\notGate[277] )) /* synthesis syn_instantiated=1, lut_function=((!D !C !B !A)+(!D !C !B A)+(!D !C B !A)+(!D !C B A)+(!D C !B !A)+(!D C !B A)+(!D C B !A)+(!D C B A)), LSE_LINE_FILE_ID=3, LSE_LCOL=13, LSE_RCOL=44, LSE_LLINE=32, LSE_RLINE=32 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(11[2:53])
    defparam I1.init = 16'b0000000011111111;
    
endmodule
//
// Verilog Description of module inverter_U803
//

module inverter_U803 (\notGate[275]_keep , \notGate[276] ) /* synthesis syn_module_defined=1 */ ;
    input \notGate[275]_keep ;
    output \notGate[276] ;
    
    wire \notGate[275]_keep  /* synthesis alspreserve=1 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(25[15:22])
    
    LUT4 I1 (.A(\notGate[275]_keep ), .B(\notGate[275]_keep ), .C(\notGate[275]_keep ), 
         .D(\notGate[275]_keep ), .Z(\notGate[276] )) /* synthesis syn_instantiated=1, lut_function=((!D !C !B !A)+(!D !C !B A)+(!D !C B !A)+(!D !C B A)+(!D C !B !A)+(!D C !B A)+(!D C B !A)+(!D C B A)), LSE_LINE_FILE_ID=3, LSE_LCOL=13, LSE_RCOL=44, LSE_LLINE=32, LSE_RLINE=32 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(11[2:53])
    defparam I1.init = 16'b0000000011111111;
    
endmodule
//
// Verilog Description of module inverter_U804
//

module inverter_U804 (\notGate[274]_keep , \notGate[275] ) /* synthesis syn_module_defined=1 */ ;
    input \notGate[274]_keep ;
    output \notGate[275] ;
    
    wire \notGate[274]_keep  /* synthesis alspreserve=1 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(25[15:22])
    
    LUT4 I1 (.A(\notGate[274]_keep ), .B(\notGate[274]_keep ), .C(\notGate[274]_keep ), 
         .D(\notGate[274]_keep ), .Z(\notGate[275] )) /* synthesis syn_instantiated=1, lut_function=((!D !C !B !A)+(!D !C !B A)+(!D !C B !A)+(!D !C B A)+(!D C !B !A)+(!D C !B A)+(!D C B !A)+(!D C B A)), LSE_LINE_FILE_ID=3, LSE_LCOL=13, LSE_RCOL=44, LSE_LLINE=32, LSE_RLINE=32 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(11[2:53])
    defparam I1.init = 16'b0000000011111111;
    
endmodule
//
// Verilog Description of module inverter_U805
//

module inverter_U805 (\notGate[273]_keep , \notGate[274] ) /* synthesis syn_module_defined=1 */ ;
    input \notGate[273]_keep ;
    output \notGate[274] ;
    
    wire \notGate[273]_keep  /* synthesis alspreserve=1 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(25[15:22])
    
    LUT4 I1 (.A(\notGate[273]_keep ), .B(\notGate[273]_keep ), .C(\notGate[273]_keep ), 
         .D(\notGate[273]_keep ), .Z(\notGate[274] )) /* synthesis syn_instantiated=1, lut_function=((!D !C !B !A)+(!D !C !B A)+(!D !C B !A)+(!D !C B A)+(!D C !B !A)+(!D C !B A)+(!D C B !A)+(!D C B A)), LSE_LINE_FILE_ID=3, LSE_LCOL=13, LSE_RCOL=44, LSE_LLINE=32, LSE_RLINE=32 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(11[2:53])
    defparam I1.init = 16'b0000000011111111;
    
endmodule
//
// Verilog Description of module inverter_U806
//

module inverter_U806 (\notGate[272]_keep , \notGate[273] ) /* synthesis syn_module_defined=1 */ ;
    input \notGate[272]_keep ;
    output \notGate[273] ;
    
    wire \notGate[272]_keep  /* synthesis alspreserve=1 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(25[15:22])
    
    LUT4 I1 (.A(\notGate[272]_keep ), .B(\notGate[272]_keep ), .C(\notGate[272]_keep ), 
         .D(\notGate[272]_keep ), .Z(\notGate[273] )) /* synthesis syn_instantiated=1, lut_function=((!D !C !B !A)+(!D !C !B A)+(!D !C B !A)+(!D !C B A)+(!D C !B !A)+(!D C !B A)+(!D C B !A)+(!D C B A)), LSE_LINE_FILE_ID=3, LSE_LCOL=13, LSE_RCOL=44, LSE_LLINE=32, LSE_RLINE=32 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(11[2:53])
    defparam I1.init = 16'b0000000011111111;
    
endmodule
//
// Verilog Description of module inverter_U807
//

module inverter_U807 (\notGate[271]_keep , \notGate[272] ) /* synthesis syn_module_defined=1 */ ;
    input \notGate[271]_keep ;
    output \notGate[272] ;
    
    wire \notGate[271]_keep  /* synthesis alspreserve=1 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(25[15:22])
    
    LUT4 I1 (.A(\notGate[271]_keep ), .B(\notGate[271]_keep ), .C(\notGate[271]_keep ), 
         .D(\notGate[271]_keep ), .Z(\notGate[272] )) /* synthesis syn_instantiated=1, lut_function=((!D !C !B !A)+(!D !C !B A)+(!D !C B !A)+(!D !C B A)+(!D C !B !A)+(!D C !B A)+(!D C B !A)+(!D C B A)), LSE_LINE_FILE_ID=3, LSE_LCOL=13, LSE_RCOL=44, LSE_LLINE=32, LSE_RLINE=32 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(11[2:53])
    defparam I1.init = 16'b0000000011111111;
    
endmodule
//
// Verilog Description of module inverter_U808
//

module inverter_U808 (\notGate[270]_keep , \notGate[271] ) /* synthesis syn_module_defined=1 */ ;
    input \notGate[270]_keep ;
    output \notGate[271] ;
    
    wire \notGate[270]_keep  /* synthesis alspreserve=1 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(25[15:22])
    
    LUT4 I1 (.A(\notGate[270]_keep ), .B(\notGate[270]_keep ), .C(\notGate[270]_keep ), 
         .D(\notGate[270]_keep ), .Z(\notGate[271] )) /* synthesis syn_instantiated=1, lut_function=((!D !C !B !A)+(!D !C !B A)+(!D !C B !A)+(!D !C B A)+(!D C !B !A)+(!D C !B A)+(!D C B !A)+(!D C B A)), LSE_LINE_FILE_ID=3, LSE_LCOL=13, LSE_RCOL=44, LSE_LLINE=32, LSE_RLINE=32 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(11[2:53])
    defparam I1.init = 16'b0000000011111111;
    
endmodule
//
// Verilog Description of module inverter_U809
//

module inverter_U809 (\notGate[269]_keep , \notGate[270] ) /* synthesis syn_module_defined=1 */ ;
    input \notGate[269]_keep ;
    output \notGate[270] ;
    
    wire \notGate[269]_keep  /* synthesis alspreserve=1 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(25[15:22])
    
    LUT4 I1 (.A(\notGate[269]_keep ), .B(\notGate[269]_keep ), .C(\notGate[269]_keep ), 
         .D(\notGate[269]_keep ), .Z(\notGate[270] )) /* synthesis syn_instantiated=1, lut_function=((!D !C !B !A)+(!D !C !B A)+(!D !C B !A)+(!D !C B A)+(!D C !B !A)+(!D C !B A)+(!D C B !A)+(!D C B A)), LSE_LINE_FILE_ID=3, LSE_LCOL=13, LSE_RCOL=44, LSE_LLINE=32, LSE_RLINE=32 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(11[2:53])
    defparam I1.init = 16'b0000000011111111;
    
endmodule
//
// Verilog Description of module inverter_U810
//

module inverter_U810 (\notGate[25]_keep , \notGate[26] ) /* synthesis syn_module_defined=1 */ ;
    input \notGate[25]_keep ;
    output \notGate[26] ;
    
    wire \notGate[25]_keep  /* synthesis alspreserve=1 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(25[15:22])
    
    LUT4 I1 (.A(\notGate[25]_keep ), .B(\notGate[25]_keep ), .C(\notGate[25]_keep ), 
         .D(\notGate[25]_keep ), .Z(\notGate[26] )) /* synthesis syn_instantiated=1, lut_function=((!D !C !B !A)+(!D !C !B A)+(!D !C B !A)+(!D !C B A)+(!D C !B !A)+(!D C !B A)+(!D C B !A)+(!D C B A)), LSE_LINE_FILE_ID=3, LSE_LCOL=13, LSE_RCOL=44, LSE_LLINE=32, LSE_RLINE=32 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(11[2:53])
    defparam I1.init = 16'b0000000011111111;
    
endmodule
//
// Verilog Description of module inverter_U811
//

module inverter_U811 (\notGate[268]_keep , \notGate[269] ) /* synthesis syn_module_defined=1 */ ;
    input \notGate[268]_keep ;
    output \notGate[269] ;
    
    wire \notGate[268]_keep  /* synthesis alspreserve=1 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(25[15:22])
    
    LUT4 I1 (.A(\notGate[268]_keep ), .B(\notGate[268]_keep ), .C(\notGate[268]_keep ), 
         .D(\notGate[268]_keep ), .Z(\notGate[269] )) /* synthesis syn_instantiated=1, lut_function=((!D !C !B !A)+(!D !C !B A)+(!D !C B !A)+(!D !C B A)+(!D C !B !A)+(!D C !B A)+(!D C B !A)+(!D C B A)), LSE_LINE_FILE_ID=3, LSE_LCOL=13, LSE_RCOL=44, LSE_LLINE=32, LSE_RLINE=32 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(11[2:53])
    defparam I1.init = 16'b0000000011111111;
    
endmodule
//
// Verilog Description of module inverter_U812
//

module inverter_U812 (\notGate[267]_keep , \notGate[268] ) /* synthesis syn_module_defined=1 */ ;
    input \notGate[267]_keep ;
    output \notGate[268] ;
    
    wire \notGate[267]_keep  /* synthesis alspreserve=1 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(25[15:22])
    
    LUT4 I1 (.A(\notGate[267]_keep ), .B(\notGate[267]_keep ), .C(\notGate[267]_keep ), 
         .D(\notGate[267]_keep ), .Z(\notGate[268] )) /* synthesis syn_instantiated=1, lut_function=((!D !C !B !A)+(!D !C !B A)+(!D !C B !A)+(!D !C B A)+(!D C !B !A)+(!D C !B A)+(!D C B !A)+(!D C B A)), LSE_LINE_FILE_ID=3, LSE_LCOL=13, LSE_RCOL=44, LSE_LLINE=32, LSE_RLINE=32 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(11[2:53])
    defparam I1.init = 16'b0000000011111111;
    
endmodule
//
// Verilog Description of module inverter_U813
//

module inverter_U813 (\notGate[266]_keep , \notGate[267] ) /* synthesis syn_module_defined=1 */ ;
    input \notGate[266]_keep ;
    output \notGate[267] ;
    
    wire \notGate[266]_keep  /* synthesis alspreserve=1 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(25[15:22])
    
    LUT4 I1 (.A(\notGate[266]_keep ), .B(\notGate[266]_keep ), .C(\notGate[266]_keep ), 
         .D(\notGate[266]_keep ), .Z(\notGate[267] )) /* synthesis syn_instantiated=1, lut_function=((!D !C !B !A)+(!D !C !B A)+(!D !C B !A)+(!D !C B A)+(!D C !B !A)+(!D C !B A)+(!D C B !A)+(!D C B A)), LSE_LINE_FILE_ID=3, LSE_LCOL=13, LSE_RCOL=44, LSE_LLINE=32, LSE_RLINE=32 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(11[2:53])
    defparam I1.init = 16'b0000000011111111;
    
endmodule
//
// Verilog Description of module inverter_U814
//

module inverter_U814 (\notGate[265]_keep , \notGate[266] ) /* synthesis syn_module_defined=1 */ ;
    input \notGate[265]_keep ;
    output \notGate[266] ;
    
    wire \notGate[265]_keep  /* synthesis alspreserve=1 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(25[15:22])
    
    LUT4 I1 (.A(\notGate[265]_keep ), .B(\notGate[265]_keep ), .C(\notGate[265]_keep ), 
         .D(\notGate[265]_keep ), .Z(\notGate[266] )) /* synthesis syn_instantiated=1, lut_function=((!D !C !B !A)+(!D !C !B A)+(!D !C B !A)+(!D !C B A)+(!D C !B !A)+(!D C !B A)+(!D C B !A)+(!D C B A)), LSE_LINE_FILE_ID=3, LSE_LCOL=13, LSE_RCOL=44, LSE_LLINE=32, LSE_RLINE=32 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(11[2:53])
    defparam I1.init = 16'b0000000011111111;
    
endmodule
//
// Verilog Description of module inverter_U815
//

module inverter_U815 (\notGate[264]_keep , \notGate[265] ) /* synthesis syn_module_defined=1 */ ;
    input \notGate[264]_keep ;
    output \notGate[265] ;
    
    wire \notGate[264]_keep  /* synthesis alspreserve=1 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(25[15:22])
    
    LUT4 I1 (.A(\notGate[264]_keep ), .B(\notGate[264]_keep ), .C(\notGate[264]_keep ), 
         .D(\notGate[264]_keep ), .Z(\notGate[265] )) /* synthesis syn_instantiated=1, lut_function=((!D !C !B !A)+(!D !C !B A)+(!D !C B !A)+(!D !C B A)+(!D C !B !A)+(!D C !B A)+(!D C B !A)+(!D C B A)), LSE_LINE_FILE_ID=3, LSE_LCOL=13, LSE_RCOL=44, LSE_LLINE=32, LSE_RLINE=32 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(11[2:53])
    defparam I1.init = 16'b0000000011111111;
    
endmodule
//
// Verilog Description of module inverter_U816
//

module inverter_U816 (\notGate[263]_keep , \notGate[264] ) /* synthesis syn_module_defined=1 */ ;
    input \notGate[263]_keep ;
    output \notGate[264] ;
    
    wire \notGate[263]_keep  /* synthesis alspreserve=1 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(25[15:22])
    
    LUT4 I1 (.A(\notGate[263]_keep ), .B(\notGate[263]_keep ), .C(\notGate[263]_keep ), 
         .D(\notGate[263]_keep ), .Z(\notGate[264] )) /* synthesis syn_instantiated=1, lut_function=((!D !C !B !A)+(!D !C !B A)+(!D !C B !A)+(!D !C B A)+(!D C !B !A)+(!D C !B A)+(!D C B !A)+(!D C B A)), LSE_LINE_FILE_ID=3, LSE_LCOL=13, LSE_RCOL=44, LSE_LLINE=32, LSE_RLINE=32 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(11[2:53])
    defparam I1.init = 16'b0000000011111111;
    
endmodule
//
// Verilog Description of module inverter_U817
//

module inverter_U817 (\notGate[262]_keep , \notGate[263] ) /* synthesis syn_module_defined=1 */ ;
    input \notGate[262]_keep ;
    output \notGate[263] ;
    
    wire \notGate[262]_keep  /* synthesis alspreserve=1 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(25[15:22])
    
    LUT4 I1 (.A(\notGate[262]_keep ), .B(\notGate[262]_keep ), .C(\notGate[262]_keep ), 
         .D(\notGate[262]_keep ), .Z(\notGate[263] )) /* synthesis syn_instantiated=1, lut_function=((!D !C !B !A)+(!D !C !B A)+(!D !C B !A)+(!D !C B A)+(!D C !B !A)+(!D C !B A)+(!D C B !A)+(!D C B A)), LSE_LINE_FILE_ID=3, LSE_LCOL=13, LSE_RCOL=44, LSE_LLINE=32, LSE_RLINE=32 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(11[2:53])
    defparam I1.init = 16'b0000000011111111;
    
endmodule
//
// Verilog Description of module inverter_U818
//

module inverter_U818 (\notGate[261]_keep , \notGate[262] ) /* synthesis syn_module_defined=1 */ ;
    input \notGate[261]_keep ;
    output \notGate[262] ;
    
    wire \notGate[261]_keep  /* synthesis alspreserve=1 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(25[15:22])
    
    LUT4 I1 (.A(\notGate[261]_keep ), .B(\notGate[261]_keep ), .C(\notGate[261]_keep ), 
         .D(\notGate[261]_keep ), .Z(\notGate[262] )) /* synthesis syn_instantiated=1, lut_function=((!D !C !B !A)+(!D !C !B A)+(!D !C B !A)+(!D !C B A)+(!D C !B !A)+(!D C !B A)+(!D C B !A)+(!D C B A)), LSE_LINE_FILE_ID=3, LSE_LCOL=13, LSE_RCOL=44, LSE_LLINE=32, LSE_RLINE=32 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(11[2:53])
    defparam I1.init = 16'b0000000011111111;
    
endmodule
//
// Verilog Description of module inverter_U819
//

module inverter_U819 (\notGate[260]_keep , \notGate[261] ) /* synthesis syn_module_defined=1 */ ;
    input \notGate[260]_keep ;
    output \notGate[261] ;
    
    wire \notGate[260]_keep  /* synthesis alspreserve=1 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(25[15:22])
    
    LUT4 I1 (.A(\notGate[260]_keep ), .B(\notGate[260]_keep ), .C(\notGate[260]_keep ), 
         .D(\notGate[260]_keep ), .Z(\notGate[261] )) /* synthesis syn_instantiated=1, lut_function=((!D !C !B !A)+(!D !C !B A)+(!D !C B !A)+(!D !C B A)+(!D C !B !A)+(!D C !B A)+(!D C B !A)+(!D C B A)), LSE_LINE_FILE_ID=3, LSE_LCOL=13, LSE_RCOL=44, LSE_LLINE=32, LSE_RLINE=32 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(11[2:53])
    defparam I1.init = 16'b0000000011111111;
    
endmodule
//
// Verilog Description of module inverter_U820
//

module inverter_U820 (\notGate[259]_keep , \notGate[260] ) /* synthesis syn_module_defined=1 */ ;
    input \notGate[259]_keep ;
    output \notGate[260] ;
    
    wire \notGate[259]_keep  /* synthesis alspreserve=1 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(25[15:22])
    
    LUT4 I1 (.A(\notGate[259]_keep ), .B(\notGate[259]_keep ), .C(\notGate[259]_keep ), 
         .D(\notGate[259]_keep ), .Z(\notGate[260] )) /* synthesis syn_instantiated=1, lut_function=((!D !C !B !A)+(!D !C !B A)+(!D !C B !A)+(!D !C B A)+(!D C !B !A)+(!D C !B A)+(!D C B !A)+(!D C B A)), LSE_LINE_FILE_ID=3, LSE_LCOL=13, LSE_RCOL=44, LSE_LLINE=32, LSE_RLINE=32 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(11[2:53])
    defparam I1.init = 16'b0000000011111111;
    
endmodule
//
// Verilog Description of module inverter_U821
//

module inverter_U821 (\notGate[24]_keep , \notGate[25] ) /* synthesis syn_module_defined=1 */ ;
    input \notGate[24]_keep ;
    output \notGate[25] ;
    
    wire \notGate[24]_keep  /* synthesis alspreserve=1 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(25[15:22])
    
    LUT4 I1 (.A(\notGate[24]_keep ), .B(\notGate[24]_keep ), .C(\notGate[24]_keep ), 
         .D(\notGate[24]_keep ), .Z(\notGate[25] )) /* synthesis syn_instantiated=1, lut_function=((!D !C !B !A)+(!D !C !B A)+(!D !C B !A)+(!D !C B A)+(!D C !B !A)+(!D C !B A)+(!D C B !A)+(!D C B A)), LSE_LINE_FILE_ID=3, LSE_LCOL=13, LSE_RCOL=44, LSE_LLINE=32, LSE_RLINE=32 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(11[2:53])
    defparam I1.init = 16'b0000000011111111;
    
endmodule
//
// Verilog Description of module inverter_U822
//

module inverter_U822 (\notGate[258]_keep , \notGate[259] ) /* synthesis syn_module_defined=1 */ ;
    input \notGate[258]_keep ;
    output \notGate[259] ;
    
    wire \notGate[258]_keep  /* synthesis alspreserve=1 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(25[15:22])
    
    LUT4 I1 (.A(\notGate[258]_keep ), .B(\notGate[258]_keep ), .C(\notGate[258]_keep ), 
         .D(\notGate[258]_keep ), .Z(\notGate[259] )) /* synthesis syn_instantiated=1, lut_function=((!D !C !B !A)+(!D !C !B A)+(!D !C B !A)+(!D !C B A)+(!D C !B !A)+(!D C !B A)+(!D C B !A)+(!D C B A)), LSE_LINE_FILE_ID=3, LSE_LCOL=13, LSE_RCOL=44, LSE_LLINE=32, LSE_RLINE=32 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(11[2:53])
    defparam I1.init = 16'b0000000011111111;
    
endmodule
//
// Verilog Description of module inverter_U823
//

module inverter_U823 (\notGate[257]_keep , \notGate[258] ) /* synthesis syn_module_defined=1 */ ;
    input \notGate[257]_keep ;
    output \notGate[258] ;
    
    wire \notGate[257]_keep  /* synthesis alspreserve=1 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(25[15:22])
    
    LUT4 I1 (.A(\notGate[257]_keep ), .B(\notGate[257]_keep ), .C(\notGate[257]_keep ), 
         .D(\notGate[257]_keep ), .Z(\notGate[258] )) /* synthesis syn_instantiated=1, lut_function=((!D !C !B !A)+(!D !C !B A)+(!D !C B !A)+(!D !C B A)+(!D C !B !A)+(!D C !B A)+(!D C B !A)+(!D C B A)), LSE_LINE_FILE_ID=3, LSE_LCOL=13, LSE_RCOL=44, LSE_LLINE=32, LSE_RLINE=32 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(11[2:53])
    defparam I1.init = 16'b0000000011111111;
    
endmodule
//
// Verilog Description of module inverter_U824
//

module inverter_U824 (\notGate[256]_keep , \notGate[257] ) /* synthesis syn_module_defined=1 */ ;
    input \notGate[256]_keep ;
    output \notGate[257] ;
    
    wire \notGate[256]_keep  /* synthesis alspreserve=1 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(25[15:22])
    
    LUT4 I1 (.A(\notGate[256]_keep ), .B(\notGate[256]_keep ), .C(\notGate[256]_keep ), 
         .D(\notGate[256]_keep ), .Z(\notGate[257] )) /* synthesis syn_instantiated=1, lut_function=((!D !C !B !A)+(!D !C !B A)+(!D !C B !A)+(!D !C B A)+(!D C !B !A)+(!D C !B A)+(!D C B !A)+(!D C B A)), LSE_LINE_FILE_ID=3, LSE_LCOL=13, LSE_RCOL=44, LSE_LLINE=32, LSE_RLINE=32 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(11[2:53])
    defparam I1.init = 16'b0000000011111111;
    
endmodule
//
// Verilog Description of module inverter_U825
//

module inverter_U825 (\notGate[255]_keep , \notGate[256] ) /* synthesis syn_module_defined=1 */ ;
    input \notGate[255]_keep ;
    output \notGate[256] ;
    
    wire \notGate[255]_keep  /* synthesis alspreserve=1 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(25[15:22])
    
    LUT4 I1 (.A(\notGate[255]_keep ), .B(\notGate[255]_keep ), .C(\notGate[255]_keep ), 
         .D(\notGate[255]_keep ), .Z(\notGate[256] )) /* synthesis syn_instantiated=1, lut_function=((!D !C !B !A)+(!D !C !B A)+(!D !C B !A)+(!D !C B A)+(!D C !B !A)+(!D C !B A)+(!D C B !A)+(!D C B A)), LSE_LINE_FILE_ID=3, LSE_LCOL=13, LSE_RCOL=44, LSE_LLINE=32, LSE_RLINE=32 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(11[2:53])
    defparam I1.init = 16'b0000000011111111;
    
endmodule
//
// Verilog Description of module inverter_U826
//

module inverter_U826 (\notGate[254]_keep , \notGate[255] ) /* synthesis syn_module_defined=1 */ ;
    input \notGate[254]_keep ;
    output \notGate[255] ;
    
    wire \notGate[254]_keep  /* synthesis alspreserve=1 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(25[15:22])
    
    LUT4 I1 (.A(\notGate[254]_keep ), .B(\notGate[254]_keep ), .C(\notGate[254]_keep ), 
         .D(\notGate[254]_keep ), .Z(\notGate[255] )) /* synthesis syn_instantiated=1, lut_function=((!D !C !B !A)+(!D !C !B A)+(!D !C B !A)+(!D !C B A)+(!D C !B !A)+(!D C !B A)+(!D C B !A)+(!D C B A)), LSE_LINE_FILE_ID=3, LSE_LCOL=13, LSE_RCOL=44, LSE_LLINE=32, LSE_RLINE=32 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(11[2:53])
    defparam I1.init = 16'b0000000011111111;
    
endmodule
//
// Verilog Description of module inverter_U827
//

module inverter_U827 (\notGate[253]_keep , \notGate[254] ) /* synthesis syn_module_defined=1 */ ;
    input \notGate[253]_keep ;
    output \notGate[254] ;
    
    wire \notGate[253]_keep  /* synthesis alspreserve=1 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(25[15:22])
    
    LUT4 I1 (.A(\notGate[253]_keep ), .B(\notGate[253]_keep ), .C(\notGate[253]_keep ), 
         .D(\notGate[253]_keep ), .Z(\notGate[254] )) /* synthesis syn_instantiated=1, lut_function=((!D !C !B !A)+(!D !C !B A)+(!D !C B !A)+(!D !C B A)+(!D C !B !A)+(!D C !B A)+(!D C B !A)+(!D C B A)), LSE_LINE_FILE_ID=3, LSE_LCOL=13, LSE_RCOL=44, LSE_LLINE=32, LSE_RLINE=32 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(11[2:53])
    defparam I1.init = 16'b0000000011111111;
    
endmodule
//
// Verilog Description of module inverter_U828
//

module inverter_U828 (\notGate[252]_keep , \notGate[253] ) /* synthesis syn_module_defined=1 */ ;
    input \notGate[252]_keep ;
    output \notGate[253] ;
    
    wire \notGate[252]_keep  /* synthesis alspreserve=1 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(25[15:22])
    
    LUT4 I1 (.A(\notGate[252]_keep ), .B(\notGate[252]_keep ), .C(\notGate[252]_keep ), 
         .D(\notGate[252]_keep ), .Z(\notGate[253] )) /* synthesis syn_instantiated=1, lut_function=((!D !C !B !A)+(!D !C !B A)+(!D !C B !A)+(!D !C B A)+(!D C !B !A)+(!D C !B A)+(!D C B !A)+(!D C B A)), LSE_LINE_FILE_ID=3, LSE_LCOL=13, LSE_RCOL=44, LSE_LLINE=32, LSE_RLINE=32 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(11[2:53])
    defparam I1.init = 16'b0000000011111111;
    
endmodule
//
// Verilog Description of module inverter_U829
//

module inverter_U829 (\notGate[251]_keep , \notGate[252] ) /* synthesis syn_module_defined=1 */ ;
    input \notGate[251]_keep ;
    output \notGate[252] ;
    
    wire \notGate[251]_keep  /* synthesis alspreserve=1 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(25[15:22])
    
    LUT4 I1 (.A(\notGate[251]_keep ), .B(\notGate[251]_keep ), .C(\notGate[251]_keep ), 
         .D(\notGate[251]_keep ), .Z(\notGate[252] )) /* synthesis syn_instantiated=1, lut_function=((!D !C !B !A)+(!D !C !B A)+(!D !C B !A)+(!D !C B A)+(!D C !B !A)+(!D C !B A)+(!D C B !A)+(!D C B A)), LSE_LINE_FILE_ID=3, LSE_LCOL=13, LSE_RCOL=44, LSE_LLINE=32, LSE_RLINE=32 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(11[2:53])
    defparam I1.init = 16'b0000000011111111;
    
endmodule
//
// Verilog Description of module inverter_U830
//

module inverter_U830 (\notGate[250]_keep , \notGate[251] ) /* synthesis syn_module_defined=1 */ ;
    input \notGate[250]_keep ;
    output \notGate[251] ;
    
    wire \notGate[250]_keep  /* synthesis alspreserve=1 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(25[15:22])
    
    LUT4 I1 (.A(\notGate[250]_keep ), .B(\notGate[250]_keep ), .C(\notGate[250]_keep ), 
         .D(\notGate[250]_keep ), .Z(\notGate[251] )) /* synthesis syn_instantiated=1, lut_function=((!D !C !B !A)+(!D !C !B A)+(!D !C B !A)+(!D !C B A)+(!D C !B !A)+(!D C !B A)+(!D C B !A)+(!D C B A)), LSE_LINE_FILE_ID=3, LSE_LCOL=13, LSE_RCOL=44, LSE_LLINE=32, LSE_RLINE=32 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(11[2:53])
    defparam I1.init = 16'b0000000011111111;
    
endmodule
//
// Verilog Description of module inverter_U831
//

module inverter_U831 (\notGate[249]_keep , \notGate[250] ) /* synthesis syn_module_defined=1 */ ;
    input \notGate[249]_keep ;
    output \notGate[250] ;
    
    wire \notGate[249]_keep  /* synthesis alspreserve=1 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(25[15:22])
    
    LUT4 I1 (.A(\notGate[249]_keep ), .B(\notGate[249]_keep ), .C(\notGate[249]_keep ), 
         .D(\notGate[249]_keep ), .Z(\notGate[250] )) /* synthesis syn_instantiated=1, lut_function=((!D !C !B !A)+(!D !C !B A)+(!D !C B !A)+(!D !C B A)+(!D C !B !A)+(!D C !B A)+(!D C B !A)+(!D C B A)), LSE_LINE_FILE_ID=3, LSE_LCOL=13, LSE_RCOL=44, LSE_LLINE=32, LSE_RLINE=32 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(11[2:53])
    defparam I1.init = 16'b0000000011111111;
    
endmodule
//
// Verilog Description of module inverter_U832
//

module inverter_U832 (\notGate[23]_keep , \notGate[24] ) /* synthesis syn_module_defined=1 */ ;
    input \notGate[23]_keep ;
    output \notGate[24] ;
    
    wire \notGate[23]_keep  /* synthesis alspreserve=1 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(25[15:22])
    
    LUT4 I1 (.A(\notGate[23]_keep ), .B(\notGate[23]_keep ), .C(\notGate[23]_keep ), 
         .D(\notGate[23]_keep ), .Z(\notGate[24] )) /* synthesis syn_instantiated=1, lut_function=((!D !C !B !A)+(!D !C !B A)+(!D !C B !A)+(!D !C B A)+(!D C !B !A)+(!D C !B A)+(!D C B !A)+(!D C B A)), LSE_LINE_FILE_ID=3, LSE_LCOL=13, LSE_RCOL=44, LSE_LLINE=32, LSE_RLINE=32 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(11[2:53])
    defparam I1.init = 16'b0000000011111111;
    
endmodule
//
// Verilog Description of module inverter_U833
//

module inverter_U833 (\notGate[248]_keep , \notGate[249] ) /* synthesis syn_module_defined=1 */ ;
    input \notGate[248]_keep ;
    output \notGate[249] ;
    
    wire \notGate[248]_keep  /* synthesis alspreserve=1 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(25[15:22])
    
    LUT4 I1 (.A(\notGate[248]_keep ), .B(\notGate[248]_keep ), .C(\notGate[248]_keep ), 
         .D(\notGate[248]_keep ), .Z(\notGate[249] )) /* synthesis syn_instantiated=1, lut_function=((!D !C !B !A)+(!D !C !B A)+(!D !C B !A)+(!D !C B A)+(!D C !B !A)+(!D C !B A)+(!D C B !A)+(!D C B A)), LSE_LINE_FILE_ID=3, LSE_LCOL=13, LSE_RCOL=44, LSE_LLINE=32, LSE_RLINE=32 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(11[2:53])
    defparam I1.init = 16'b0000000011111111;
    
endmodule
//
// Verilog Description of module inverter_U834
//

module inverter_U834 (\notGate[247]_keep , \notGate[248] ) /* synthesis syn_module_defined=1 */ ;
    input \notGate[247]_keep ;
    output \notGate[248] ;
    
    wire \notGate[247]_keep  /* synthesis alspreserve=1 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(25[15:22])
    
    LUT4 I1 (.A(\notGate[247]_keep ), .B(\notGate[247]_keep ), .C(\notGate[247]_keep ), 
         .D(\notGate[247]_keep ), .Z(\notGate[248] )) /* synthesis syn_instantiated=1, lut_function=((!D !C !B !A)+(!D !C !B A)+(!D !C B !A)+(!D !C B A)+(!D C !B !A)+(!D C !B A)+(!D C B !A)+(!D C B A)), LSE_LINE_FILE_ID=3, LSE_LCOL=13, LSE_RCOL=44, LSE_LLINE=32, LSE_RLINE=32 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(11[2:53])
    defparam I1.init = 16'b0000000011111111;
    
endmodule
//
// Verilog Description of module inverter_U835
//

module inverter_U835 (\notGate[246]_keep , \notGate[247] ) /* synthesis syn_module_defined=1 */ ;
    input \notGate[246]_keep ;
    output \notGate[247] ;
    
    wire \notGate[246]_keep  /* synthesis alspreserve=1 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(25[15:22])
    
    LUT4 I1 (.A(\notGate[246]_keep ), .B(\notGate[246]_keep ), .C(\notGate[246]_keep ), 
         .D(\notGate[246]_keep ), .Z(\notGate[247] )) /* synthesis syn_instantiated=1, lut_function=((!D !C !B !A)+(!D !C !B A)+(!D !C B !A)+(!D !C B A)+(!D C !B !A)+(!D C !B A)+(!D C B !A)+(!D C B A)), LSE_LINE_FILE_ID=3, LSE_LCOL=13, LSE_RCOL=44, LSE_LLINE=32, LSE_RLINE=32 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(11[2:53])
    defparam I1.init = 16'b0000000011111111;
    
endmodule
//
// Verilog Description of module inverter_U836
//

module inverter_U836 (\notGate[245]_keep , \notGate[246] ) /* synthesis syn_module_defined=1 */ ;
    input \notGate[245]_keep ;
    output \notGate[246] ;
    
    wire \notGate[245]_keep  /* synthesis alspreserve=1 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(25[15:22])
    
    LUT4 I1 (.A(\notGate[245]_keep ), .B(\notGate[245]_keep ), .C(\notGate[245]_keep ), 
         .D(\notGate[245]_keep ), .Z(\notGate[246] )) /* synthesis syn_instantiated=1, lut_function=((!D !C !B !A)+(!D !C !B A)+(!D !C B !A)+(!D !C B A)+(!D C !B !A)+(!D C !B A)+(!D C B !A)+(!D C B A)), LSE_LINE_FILE_ID=3, LSE_LCOL=13, LSE_RCOL=44, LSE_LLINE=32, LSE_RLINE=32 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(11[2:53])
    defparam I1.init = 16'b0000000011111111;
    
endmodule
//
// Verilog Description of module inverter_U837
//

module inverter_U837 (\notGate[244]_keep , \notGate[245] ) /* synthesis syn_module_defined=1 */ ;
    input \notGate[244]_keep ;
    output \notGate[245] ;
    
    wire \notGate[244]_keep  /* synthesis alspreserve=1 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(25[15:22])
    
    LUT4 I1 (.A(\notGate[244]_keep ), .B(\notGate[244]_keep ), .C(\notGate[244]_keep ), 
         .D(\notGate[244]_keep ), .Z(\notGate[245] )) /* synthesis syn_instantiated=1, lut_function=((!D !C !B !A)+(!D !C !B A)+(!D !C B !A)+(!D !C B A)+(!D C !B !A)+(!D C !B A)+(!D C B !A)+(!D C B A)), LSE_LINE_FILE_ID=3, LSE_LCOL=13, LSE_RCOL=44, LSE_LLINE=32, LSE_RLINE=32 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(11[2:53])
    defparam I1.init = 16'b0000000011111111;
    
endmodule
//
// Verilog Description of module inverter_U838
//

module inverter_U838 (\notGate[243]_keep , \notGate[244] ) /* synthesis syn_module_defined=1 */ ;
    input \notGate[243]_keep ;
    output \notGate[244] ;
    
    wire \notGate[243]_keep  /* synthesis alspreserve=1 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(25[15:22])
    
    LUT4 I1 (.A(\notGate[243]_keep ), .B(\notGate[243]_keep ), .C(\notGate[243]_keep ), 
         .D(\notGate[243]_keep ), .Z(\notGate[244] )) /* synthesis syn_instantiated=1, lut_function=((!D !C !B !A)+(!D !C !B A)+(!D !C B !A)+(!D !C B A)+(!D C !B !A)+(!D C !B A)+(!D C B !A)+(!D C B A)), LSE_LINE_FILE_ID=3, LSE_LCOL=13, LSE_RCOL=44, LSE_LLINE=32, LSE_RLINE=32 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(11[2:53])
    defparam I1.init = 16'b0000000011111111;
    
endmodule
//
// Verilog Description of module inverter_U839
//

module inverter_U839 (\notGate[242]_keep , \notGate[243] ) /* synthesis syn_module_defined=1 */ ;
    input \notGate[242]_keep ;
    output \notGate[243] ;
    
    wire \notGate[242]_keep  /* synthesis alspreserve=1 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(25[15:22])
    
    LUT4 I1 (.A(\notGate[242]_keep ), .B(\notGate[242]_keep ), .C(\notGate[242]_keep ), 
         .D(\notGate[242]_keep ), .Z(\notGate[243] )) /* synthesis syn_instantiated=1, lut_function=((!D !C !B !A)+(!D !C !B A)+(!D !C B !A)+(!D !C B A)+(!D C !B !A)+(!D C !B A)+(!D C B !A)+(!D C B A)), LSE_LINE_FILE_ID=3, LSE_LCOL=13, LSE_RCOL=44, LSE_LLINE=32, LSE_RLINE=32 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(11[2:53])
    defparam I1.init = 16'b0000000011111111;
    
endmodule
//
// Verilog Description of module inverter_U840
//

module inverter_U840 (\notGate[241]_keep , \notGate[242] ) /* synthesis syn_module_defined=1 */ ;
    input \notGate[241]_keep ;
    output \notGate[242] ;
    
    wire \notGate[241]_keep  /* synthesis alspreserve=1 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(25[15:22])
    
    LUT4 I1 (.A(\notGate[241]_keep ), .B(\notGate[241]_keep ), .C(\notGate[241]_keep ), 
         .D(\notGate[241]_keep ), .Z(\notGate[242] )) /* synthesis syn_instantiated=1, lut_function=((!D !C !B !A)+(!D !C !B A)+(!D !C B !A)+(!D !C B A)+(!D C !B !A)+(!D C !B A)+(!D C B !A)+(!D C B A)), LSE_LINE_FILE_ID=3, LSE_LCOL=13, LSE_RCOL=44, LSE_LLINE=32, LSE_RLINE=32 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(11[2:53])
    defparam I1.init = 16'b0000000011111111;
    
endmodule
//
// Verilog Description of module inverter_U841
//

module inverter_U841 (\notGate[240]_keep , \notGate[241] ) /* synthesis syn_module_defined=1 */ ;
    input \notGate[240]_keep ;
    output \notGate[241] ;
    
    wire \notGate[240]_keep  /* synthesis alspreserve=1 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(25[15:22])
    
    LUT4 I1 (.A(\notGate[240]_keep ), .B(\notGate[240]_keep ), .C(\notGate[240]_keep ), 
         .D(\notGate[240]_keep ), .Z(\notGate[241] )) /* synthesis syn_instantiated=1, lut_function=((!D !C !B !A)+(!D !C !B A)+(!D !C B !A)+(!D !C B A)+(!D C !B !A)+(!D C !B A)+(!D C B !A)+(!D C B A)), LSE_LINE_FILE_ID=3, LSE_LCOL=13, LSE_RCOL=44, LSE_LLINE=32, LSE_RLINE=32 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(11[2:53])
    defparam I1.init = 16'b0000000011111111;
    
endmodule
//
// Verilog Description of module inverter_U842
//

module inverter_U842 (\notGate[239]_keep , \notGate[240] ) /* synthesis syn_module_defined=1 */ ;
    input \notGate[239]_keep ;
    output \notGate[240] ;
    
    wire \notGate[239]_keep  /* synthesis alspreserve=1 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(25[15:22])
    
    LUT4 I1 (.A(\notGate[239]_keep ), .B(\notGate[239]_keep ), .C(\notGate[239]_keep ), 
         .D(\notGate[239]_keep ), .Z(\notGate[240] )) /* synthesis syn_instantiated=1, lut_function=((!D !C !B !A)+(!D !C !B A)+(!D !C B !A)+(!D !C B A)+(!D C !B !A)+(!D C !B A)+(!D C B !A)+(!D C B A)), LSE_LINE_FILE_ID=3, LSE_LCOL=13, LSE_RCOL=44, LSE_LLINE=32, LSE_RLINE=32 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(11[2:53])
    defparam I1.init = 16'b0000000011111111;
    
endmodule
//
// Verilog Description of module inverter_U843
//

module inverter_U843 (\notGate[22]_keep , \notGate[23] ) /* synthesis syn_module_defined=1 */ ;
    input \notGate[22]_keep ;
    output \notGate[23] ;
    
    wire \notGate[22]_keep  /* synthesis alspreserve=1 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(25[15:22])
    
    LUT4 I1 (.A(\notGate[22]_keep ), .B(\notGate[22]_keep ), .C(\notGate[22]_keep ), 
         .D(\notGate[22]_keep ), .Z(\notGate[23] )) /* synthesis syn_instantiated=1, lut_function=((!D !C !B !A)+(!D !C !B A)+(!D !C B !A)+(!D !C B A)+(!D C !B !A)+(!D C !B A)+(!D C B !A)+(!D C B A)), LSE_LINE_FILE_ID=3, LSE_LCOL=13, LSE_RCOL=44, LSE_LLINE=32, LSE_RLINE=32 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(11[2:53])
    defparam I1.init = 16'b0000000011111111;
    
endmodule
//
// Verilog Description of module inverter_U844
//

module inverter_U844 (\notGate[238]_keep , \notGate[239] ) /* synthesis syn_module_defined=1 */ ;
    input \notGate[238]_keep ;
    output \notGate[239] ;
    
    wire \notGate[238]_keep  /* synthesis alspreserve=1 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(25[15:22])
    
    LUT4 I1 (.A(\notGate[238]_keep ), .B(\notGate[238]_keep ), .C(\notGate[238]_keep ), 
         .D(\notGate[238]_keep ), .Z(\notGate[239] )) /* synthesis syn_instantiated=1, lut_function=((!D !C !B !A)+(!D !C !B A)+(!D !C B !A)+(!D !C B A)+(!D C !B !A)+(!D C !B A)+(!D C B !A)+(!D C B A)), LSE_LINE_FILE_ID=3, LSE_LCOL=13, LSE_RCOL=44, LSE_LLINE=32, LSE_RLINE=32 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(11[2:53])
    defparam I1.init = 16'b0000000011111111;
    
endmodule
//
// Verilog Description of module inverter_U845
//

module inverter_U845 (\notGate[237]_keep , \notGate[238] ) /* synthesis syn_module_defined=1 */ ;
    input \notGate[237]_keep ;
    output \notGate[238] ;
    
    wire \notGate[237]_keep  /* synthesis alspreserve=1 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(25[15:22])
    
    LUT4 I1 (.A(\notGate[237]_keep ), .B(\notGate[237]_keep ), .C(\notGate[237]_keep ), 
         .D(\notGate[237]_keep ), .Z(\notGate[238] )) /* synthesis syn_instantiated=1, lut_function=((!D !C !B !A)+(!D !C !B A)+(!D !C B !A)+(!D !C B A)+(!D C !B !A)+(!D C !B A)+(!D C B !A)+(!D C B A)), LSE_LINE_FILE_ID=3, LSE_LCOL=13, LSE_RCOL=44, LSE_LLINE=32, LSE_RLINE=32 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(11[2:53])
    defparam I1.init = 16'b0000000011111111;
    
endmodule
//
// Verilog Description of module inverter_U846
//

module inverter_U846 (\notGate[236]_keep , \notGate[237] ) /* synthesis syn_module_defined=1 */ ;
    input \notGate[236]_keep ;
    output \notGate[237] ;
    
    wire \notGate[236]_keep  /* synthesis alspreserve=1 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(25[15:22])
    
    LUT4 I1 (.A(\notGate[236]_keep ), .B(\notGate[236]_keep ), .C(\notGate[236]_keep ), 
         .D(\notGate[236]_keep ), .Z(\notGate[237] )) /* synthesis syn_instantiated=1, lut_function=((!D !C !B !A)+(!D !C !B A)+(!D !C B !A)+(!D !C B A)+(!D C !B !A)+(!D C !B A)+(!D C B !A)+(!D C B A)), LSE_LINE_FILE_ID=3, LSE_LCOL=13, LSE_RCOL=44, LSE_LLINE=32, LSE_RLINE=32 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(11[2:53])
    defparam I1.init = 16'b0000000011111111;
    
endmodule
//
// Verilog Description of module inverter_U847
//

module inverter_U847 (\notGate[235]_keep , \notGate[236] ) /* synthesis syn_module_defined=1 */ ;
    input \notGate[235]_keep ;
    output \notGate[236] ;
    
    wire \notGate[235]_keep  /* synthesis alspreserve=1 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(25[15:22])
    
    LUT4 I1 (.A(\notGate[235]_keep ), .B(\notGate[235]_keep ), .C(\notGate[235]_keep ), 
         .D(\notGate[235]_keep ), .Z(\notGate[236] )) /* synthesis syn_instantiated=1, lut_function=((!D !C !B !A)+(!D !C !B A)+(!D !C B !A)+(!D !C B A)+(!D C !B !A)+(!D C !B A)+(!D C B !A)+(!D C B A)), LSE_LINE_FILE_ID=3, LSE_LCOL=13, LSE_RCOL=44, LSE_LLINE=32, LSE_RLINE=32 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(11[2:53])
    defparam I1.init = 16'b0000000011111111;
    
endmodule
//
// Verilog Description of module inverter_U848
//

module inverter_U848 (\notGate[234]_keep , \notGate[235] ) /* synthesis syn_module_defined=1 */ ;
    input \notGate[234]_keep ;
    output \notGate[235] ;
    
    wire \notGate[234]_keep  /* synthesis alspreserve=1 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(25[15:22])
    
    LUT4 I1 (.A(\notGate[234]_keep ), .B(\notGate[234]_keep ), .C(\notGate[234]_keep ), 
         .D(\notGate[234]_keep ), .Z(\notGate[235] )) /* synthesis syn_instantiated=1, lut_function=((!D !C !B !A)+(!D !C !B A)+(!D !C B !A)+(!D !C B A)+(!D C !B !A)+(!D C !B A)+(!D C B !A)+(!D C B A)), LSE_LINE_FILE_ID=3, LSE_LCOL=13, LSE_RCOL=44, LSE_LLINE=32, LSE_RLINE=32 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(11[2:53])
    defparam I1.init = 16'b0000000011111111;
    
endmodule
//
// Verilog Description of module inverter_U849
//

module inverter_U849 (\notGate[233]_keep , \notGate[234] ) /* synthesis syn_module_defined=1 */ ;
    input \notGate[233]_keep ;
    output \notGate[234] ;
    
    wire \notGate[233]_keep  /* synthesis alspreserve=1 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(25[15:22])
    
    LUT4 I1 (.A(\notGate[233]_keep ), .B(\notGate[233]_keep ), .C(\notGate[233]_keep ), 
         .D(\notGate[233]_keep ), .Z(\notGate[234] )) /* synthesis syn_instantiated=1, lut_function=((!D !C !B !A)+(!D !C !B A)+(!D !C B !A)+(!D !C B A)+(!D C !B !A)+(!D C !B A)+(!D C B !A)+(!D C B A)), LSE_LINE_FILE_ID=3, LSE_LCOL=13, LSE_RCOL=44, LSE_LLINE=32, LSE_RLINE=32 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(11[2:53])
    defparam I1.init = 16'b0000000011111111;
    
endmodule
//
// Verilog Description of module inverter_U850
//

module inverter_U850 (\notGate[232]_keep , \notGate[233] ) /* synthesis syn_module_defined=1 */ ;
    input \notGate[232]_keep ;
    output \notGate[233] ;
    
    wire \notGate[232]_keep  /* synthesis alspreserve=1 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(25[15:22])
    
    LUT4 I1 (.A(\notGate[232]_keep ), .B(\notGate[232]_keep ), .C(\notGate[232]_keep ), 
         .D(\notGate[232]_keep ), .Z(\notGate[233] )) /* synthesis syn_instantiated=1, lut_function=((!D !C !B !A)+(!D !C !B A)+(!D !C B !A)+(!D !C B A)+(!D C !B !A)+(!D C !B A)+(!D C B !A)+(!D C B A)), LSE_LINE_FILE_ID=3, LSE_LCOL=13, LSE_RCOL=44, LSE_LLINE=32, LSE_RLINE=32 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(11[2:53])
    defparam I1.init = 16'b0000000011111111;
    
endmodule
//
// Verilog Description of module inverter_U851
//

module inverter_U851 (\notGate[231]_keep , \notGate[232] ) /* synthesis syn_module_defined=1 */ ;
    input \notGate[231]_keep ;
    output \notGate[232] ;
    
    wire \notGate[231]_keep  /* synthesis alspreserve=1 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(25[15:22])
    
    LUT4 I1 (.A(\notGate[231]_keep ), .B(\notGate[231]_keep ), .C(\notGate[231]_keep ), 
         .D(\notGate[231]_keep ), .Z(\notGate[232] )) /* synthesis syn_instantiated=1, lut_function=((!D !C !B !A)+(!D !C !B A)+(!D !C B !A)+(!D !C B A)+(!D C !B !A)+(!D C !B A)+(!D C B !A)+(!D C B A)), LSE_LINE_FILE_ID=3, LSE_LCOL=13, LSE_RCOL=44, LSE_LLINE=32, LSE_RLINE=32 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(11[2:53])
    defparam I1.init = 16'b0000000011111111;
    
endmodule
//
// Verilog Description of module inverter_U852
//

module inverter_U852 (\notGate[230]_keep , \notGate[231] ) /* synthesis syn_module_defined=1 */ ;
    input \notGate[230]_keep ;
    output \notGate[231] ;
    
    wire \notGate[230]_keep  /* synthesis alspreserve=1 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(25[15:22])
    
    LUT4 I1 (.A(\notGate[230]_keep ), .B(\notGate[230]_keep ), .C(\notGate[230]_keep ), 
         .D(\notGate[230]_keep ), .Z(\notGate[231] )) /* synthesis syn_instantiated=1, lut_function=((!D !C !B !A)+(!D !C !B A)+(!D !C B !A)+(!D !C B A)+(!D C !B !A)+(!D C !B A)+(!D C B !A)+(!D C B A)), LSE_LINE_FILE_ID=3, LSE_LCOL=13, LSE_RCOL=44, LSE_LLINE=32, LSE_RLINE=32 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(11[2:53])
    defparam I1.init = 16'b0000000011111111;
    
endmodule
//
// Verilog Description of module inverter_U853
//

module inverter_U853 (\notGate[229]_keep , \notGate[230] ) /* synthesis syn_module_defined=1 */ ;
    input \notGate[229]_keep ;
    output \notGate[230] ;
    
    wire \notGate[229]_keep  /* synthesis alspreserve=1 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(25[15:22])
    
    LUT4 I1 (.A(\notGate[229]_keep ), .B(\notGate[229]_keep ), .C(\notGate[229]_keep ), 
         .D(\notGate[229]_keep ), .Z(\notGate[230] )) /* synthesis syn_instantiated=1, lut_function=((!D !C !B !A)+(!D !C !B A)+(!D !C B !A)+(!D !C B A)+(!D C !B !A)+(!D C !B A)+(!D C B !A)+(!D C B A)), LSE_LINE_FILE_ID=3, LSE_LCOL=13, LSE_RCOL=44, LSE_LLINE=32, LSE_RLINE=32 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(11[2:53])
    defparam I1.init = 16'b0000000011111111;
    
endmodule
//
// Verilog Description of module inverter_U854
//

module inverter_U854 (\notGate[21]_keep , \notGate[22] ) /* synthesis syn_module_defined=1 */ ;
    input \notGate[21]_keep ;
    output \notGate[22] ;
    
    wire \notGate[21]_keep  /* synthesis alspreserve=1 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(25[15:22])
    
    LUT4 I1 (.A(\notGate[21]_keep ), .B(\notGate[21]_keep ), .C(\notGate[21]_keep ), 
         .D(\notGate[21]_keep ), .Z(\notGate[22] )) /* synthesis syn_instantiated=1, lut_function=((!D !C !B !A)+(!D !C !B A)+(!D !C B !A)+(!D !C B A)+(!D C !B !A)+(!D C !B A)+(!D C B !A)+(!D C B A)), LSE_LINE_FILE_ID=3, LSE_LCOL=13, LSE_RCOL=44, LSE_LLINE=32, LSE_RLINE=32 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(11[2:53])
    defparam I1.init = 16'b0000000011111111;
    
endmodule
//
// Verilog Description of module inverter_U855
//

module inverter_U855 (\notGate[228]_keep , \notGate[229] ) /* synthesis syn_module_defined=1 */ ;
    input \notGate[228]_keep ;
    output \notGate[229] ;
    
    wire \notGate[228]_keep  /* synthesis alspreserve=1 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(25[15:22])
    
    LUT4 I1 (.A(\notGate[228]_keep ), .B(\notGate[228]_keep ), .C(\notGate[228]_keep ), 
         .D(\notGate[228]_keep ), .Z(\notGate[229] )) /* synthesis syn_instantiated=1, lut_function=((!D !C !B !A)+(!D !C !B A)+(!D !C B !A)+(!D !C B A)+(!D C !B !A)+(!D C !B A)+(!D C B !A)+(!D C B A)), LSE_LINE_FILE_ID=3, LSE_LCOL=13, LSE_RCOL=44, LSE_LLINE=32, LSE_RLINE=32 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(11[2:53])
    defparam I1.init = 16'b0000000011111111;
    
endmodule
//
// Verilog Description of module inverter_U856
//

module inverter_U856 (\notGate[227]_keep , \notGate[228] ) /* synthesis syn_module_defined=1 */ ;
    input \notGate[227]_keep ;
    output \notGate[228] ;
    
    wire \notGate[227]_keep  /* synthesis alspreserve=1 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(25[15:22])
    
    LUT4 I1 (.A(\notGate[227]_keep ), .B(\notGate[227]_keep ), .C(\notGate[227]_keep ), 
         .D(\notGate[227]_keep ), .Z(\notGate[228] )) /* synthesis syn_instantiated=1, lut_function=((!D !C !B !A)+(!D !C !B A)+(!D !C B !A)+(!D !C B A)+(!D C !B !A)+(!D C !B A)+(!D C B !A)+(!D C B A)), LSE_LINE_FILE_ID=3, LSE_LCOL=13, LSE_RCOL=44, LSE_LLINE=32, LSE_RLINE=32 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(11[2:53])
    defparam I1.init = 16'b0000000011111111;
    
endmodule
//
// Verilog Description of module inverter_U857
//

module inverter_U857 (\notGate[226]_keep , \notGate[227] ) /* synthesis syn_module_defined=1 */ ;
    input \notGate[226]_keep ;
    output \notGate[227] ;
    
    wire \notGate[226]_keep  /* synthesis alspreserve=1 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(25[15:22])
    
    LUT4 I1 (.A(\notGate[226]_keep ), .B(\notGate[226]_keep ), .C(\notGate[226]_keep ), 
         .D(\notGate[226]_keep ), .Z(\notGate[227] )) /* synthesis syn_instantiated=1, lut_function=((!D !C !B !A)+(!D !C !B A)+(!D !C B !A)+(!D !C B A)+(!D C !B !A)+(!D C !B A)+(!D C B !A)+(!D C B A)), LSE_LINE_FILE_ID=3, LSE_LCOL=13, LSE_RCOL=44, LSE_LLINE=32, LSE_RLINE=32 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(11[2:53])
    defparam I1.init = 16'b0000000011111111;
    
endmodule
//
// Verilog Description of module inverter_U858
//

module inverter_U858 (\notGate[225]_keep , \notGate[226] ) /* synthesis syn_module_defined=1 */ ;
    input \notGate[225]_keep ;
    output \notGate[226] ;
    
    wire \notGate[225]_keep  /* synthesis alspreserve=1 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(25[15:22])
    
    LUT4 I1 (.A(\notGate[225]_keep ), .B(\notGate[225]_keep ), .C(\notGate[225]_keep ), 
         .D(\notGate[225]_keep ), .Z(\notGate[226] )) /* synthesis syn_instantiated=1, lut_function=((!D !C !B !A)+(!D !C !B A)+(!D !C B !A)+(!D !C B A)+(!D C !B !A)+(!D C !B A)+(!D C B !A)+(!D C B A)), LSE_LINE_FILE_ID=3, LSE_LCOL=13, LSE_RCOL=44, LSE_LLINE=32, LSE_RLINE=32 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(11[2:53])
    defparam I1.init = 16'b0000000011111111;
    
endmodule
//
// Verilog Description of module inverter_U859
//

module inverter_U859 (\notGate[224]_keep , \notGate[225] ) /* synthesis syn_module_defined=1 */ ;
    input \notGate[224]_keep ;
    output \notGate[225] ;
    
    wire \notGate[224]_keep  /* synthesis alspreserve=1 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(25[15:22])
    
    LUT4 I1 (.A(\notGate[224]_keep ), .B(\notGate[224]_keep ), .C(\notGate[224]_keep ), 
         .D(\notGate[224]_keep ), .Z(\notGate[225] )) /* synthesis syn_instantiated=1, lut_function=((!D !C !B !A)+(!D !C !B A)+(!D !C B !A)+(!D !C B A)+(!D C !B !A)+(!D C !B A)+(!D C B !A)+(!D C B A)), LSE_LINE_FILE_ID=3, LSE_LCOL=13, LSE_RCOL=44, LSE_LLINE=32, LSE_RLINE=32 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(11[2:53])
    defparam I1.init = 16'b0000000011111111;
    
endmodule
//
// Verilog Description of module inverter_U860
//

module inverter_U860 (\notGate[223]_keep , \notGate[224] ) /* synthesis syn_module_defined=1 */ ;
    input \notGate[223]_keep ;
    output \notGate[224] ;
    
    wire \notGate[223]_keep  /* synthesis alspreserve=1 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(25[15:22])
    
    LUT4 I1 (.A(\notGate[223]_keep ), .B(\notGate[223]_keep ), .C(\notGate[223]_keep ), 
         .D(\notGate[223]_keep ), .Z(\notGate[224] )) /* synthesis syn_instantiated=1, lut_function=((!D !C !B !A)+(!D !C !B A)+(!D !C B !A)+(!D !C B A)+(!D C !B !A)+(!D C !B A)+(!D C B !A)+(!D C B A)), LSE_LINE_FILE_ID=3, LSE_LCOL=13, LSE_RCOL=44, LSE_LLINE=32, LSE_RLINE=32 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(11[2:53])
    defparam I1.init = 16'b0000000011111111;
    
endmodule
//
// Verilog Description of module inverter_U861
//

module inverter_U861 (\notGate[222]_keep , \notGate[223] ) /* synthesis syn_module_defined=1 */ ;
    input \notGate[222]_keep ;
    output \notGate[223] ;
    
    wire \notGate[222]_keep  /* synthesis alspreserve=1 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(25[15:22])
    
    LUT4 I1 (.A(\notGate[222]_keep ), .B(\notGate[222]_keep ), .C(\notGate[222]_keep ), 
         .D(\notGate[222]_keep ), .Z(\notGate[223] )) /* synthesis syn_instantiated=1, lut_function=((!D !C !B !A)+(!D !C !B A)+(!D !C B !A)+(!D !C B A)+(!D C !B !A)+(!D C !B A)+(!D C B !A)+(!D C B A)), LSE_LINE_FILE_ID=3, LSE_LCOL=13, LSE_RCOL=44, LSE_LLINE=32, LSE_RLINE=32 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(11[2:53])
    defparam I1.init = 16'b0000000011111111;
    
endmodule
//
// Verilog Description of module inverter_U862
//

module inverter_U862 (\notGate[221]_keep , \notGate[222] ) /* synthesis syn_module_defined=1 */ ;
    input \notGate[221]_keep ;
    output \notGate[222] ;
    
    wire \notGate[221]_keep  /* synthesis alspreserve=1 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(25[15:22])
    
    LUT4 I1 (.A(\notGate[221]_keep ), .B(\notGate[221]_keep ), .C(\notGate[221]_keep ), 
         .D(\notGate[221]_keep ), .Z(\notGate[222] )) /* synthesis syn_instantiated=1, lut_function=((!D !C !B !A)+(!D !C !B A)+(!D !C B !A)+(!D !C B A)+(!D C !B !A)+(!D C !B A)+(!D C B !A)+(!D C B A)), LSE_LINE_FILE_ID=3, LSE_LCOL=13, LSE_RCOL=44, LSE_LLINE=32, LSE_RLINE=32 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(11[2:53])
    defparam I1.init = 16'b0000000011111111;
    
endmodule
//
// Verilog Description of module inverter_U863
//

module inverter_U863 (\notGate[220]_keep , \notGate[221] ) /* synthesis syn_module_defined=1 */ ;
    input \notGate[220]_keep ;
    output \notGate[221] ;
    
    wire \notGate[220]_keep  /* synthesis alspreserve=1 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(25[15:22])
    
    LUT4 I1 (.A(\notGate[220]_keep ), .B(\notGate[220]_keep ), .C(\notGate[220]_keep ), 
         .D(\notGate[220]_keep ), .Z(\notGate[221] )) /* synthesis syn_instantiated=1, lut_function=((!D !C !B !A)+(!D !C !B A)+(!D !C B !A)+(!D !C B A)+(!D C !B !A)+(!D C !B A)+(!D C B !A)+(!D C B A)), LSE_LINE_FILE_ID=3, LSE_LCOL=13, LSE_RCOL=44, LSE_LLINE=32, LSE_RLINE=32 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(11[2:53])
    defparam I1.init = 16'b0000000011111111;
    
endmodule
//
// Verilog Description of module inverter_U864
//

module inverter_U864 (\notGate[219]_keep , \notGate[220] ) /* synthesis syn_module_defined=1 */ ;
    input \notGate[219]_keep ;
    output \notGate[220] ;
    
    wire \notGate[219]_keep  /* synthesis alspreserve=1 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(25[15:22])
    
    LUT4 I1 (.A(\notGate[219]_keep ), .B(\notGate[219]_keep ), .C(\notGate[219]_keep ), 
         .D(\notGate[219]_keep ), .Z(\notGate[220] )) /* synthesis syn_instantiated=1, lut_function=((!D !C !B !A)+(!D !C !B A)+(!D !C B !A)+(!D !C B A)+(!D C !B !A)+(!D C !B A)+(!D C B !A)+(!D C B A)), LSE_LINE_FILE_ID=3, LSE_LCOL=13, LSE_RCOL=44, LSE_LLINE=32, LSE_RLINE=32 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(11[2:53])
    defparam I1.init = 16'b0000000011111111;
    
endmodule
//
// Verilog Description of module inverter_U865
//

module inverter_U865 (\notGate[20]_keep , \notGate[21] ) /* synthesis syn_module_defined=1 */ ;
    input \notGate[20]_keep ;
    output \notGate[21] ;
    
    wire \notGate[20]_keep  /* synthesis alspreserve=1 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(25[15:22])
    
    LUT4 I1 (.A(\notGate[20]_keep ), .B(\notGate[20]_keep ), .C(\notGate[20]_keep ), 
         .D(\notGate[20]_keep ), .Z(\notGate[21] )) /* synthesis syn_instantiated=1, lut_function=((!D !C !B !A)+(!D !C !B A)+(!D !C B !A)+(!D !C B A)+(!D C !B !A)+(!D C !B A)+(!D C B !A)+(!D C B A)), LSE_LINE_FILE_ID=3, LSE_LCOL=13, LSE_RCOL=44, LSE_LLINE=32, LSE_RLINE=32 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(11[2:53])
    defparam I1.init = 16'b0000000011111111;
    
endmodule
//
// Verilog Description of module inverter_U866
//

module inverter_U866 (\notGate[218]_keep , \notGate[219] ) /* synthesis syn_module_defined=1 */ ;
    input \notGate[218]_keep ;
    output \notGate[219] ;
    
    wire \notGate[218]_keep  /* synthesis alspreserve=1 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(25[15:22])
    
    LUT4 I1 (.A(\notGate[218]_keep ), .B(\notGate[218]_keep ), .C(\notGate[218]_keep ), 
         .D(\notGate[218]_keep ), .Z(\notGate[219] )) /* synthesis syn_instantiated=1, lut_function=((!D !C !B !A)+(!D !C !B A)+(!D !C B !A)+(!D !C B A)+(!D C !B !A)+(!D C !B A)+(!D C B !A)+(!D C B A)), LSE_LINE_FILE_ID=3, LSE_LCOL=13, LSE_RCOL=44, LSE_LLINE=32, LSE_RLINE=32 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(11[2:53])
    defparam I1.init = 16'b0000000011111111;
    
endmodule
//
// Verilog Description of module inverter_U867
//

module inverter_U867 (\notGate[217]_keep , \notGate[218] ) /* synthesis syn_module_defined=1 */ ;
    input \notGate[217]_keep ;
    output \notGate[218] ;
    
    wire \notGate[217]_keep  /* synthesis alspreserve=1 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(25[15:22])
    
    LUT4 I1 (.A(\notGate[217]_keep ), .B(\notGate[217]_keep ), .C(\notGate[217]_keep ), 
         .D(\notGate[217]_keep ), .Z(\notGate[218] )) /* synthesis syn_instantiated=1, lut_function=((!D !C !B !A)+(!D !C !B A)+(!D !C B !A)+(!D !C B A)+(!D C !B !A)+(!D C !B A)+(!D C B !A)+(!D C B A)), LSE_LINE_FILE_ID=3, LSE_LCOL=13, LSE_RCOL=44, LSE_LLINE=32, LSE_RLINE=32 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(11[2:53])
    defparam I1.init = 16'b0000000011111111;
    
endmodule
//
// Verilog Description of module inverter_U868
//

module inverter_U868 (\notGate[216]_keep , \notGate[217] ) /* synthesis syn_module_defined=1 */ ;
    input \notGate[216]_keep ;
    output \notGate[217] ;
    
    wire \notGate[216]_keep  /* synthesis alspreserve=1 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(25[15:22])
    
    LUT4 I1 (.A(\notGate[216]_keep ), .B(\notGate[216]_keep ), .C(\notGate[216]_keep ), 
         .D(\notGate[216]_keep ), .Z(\notGate[217] )) /* synthesis syn_instantiated=1, lut_function=((!D !C !B !A)+(!D !C !B A)+(!D !C B !A)+(!D !C B A)+(!D C !B !A)+(!D C !B A)+(!D C B !A)+(!D C B A)), LSE_LINE_FILE_ID=3, LSE_LCOL=13, LSE_RCOL=44, LSE_LLINE=32, LSE_RLINE=32 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(11[2:53])
    defparam I1.init = 16'b0000000011111111;
    
endmodule
//
// Verilog Description of module inverter_U869
//

module inverter_U869 (\notGate[215]_keep , \notGate[216] ) /* synthesis syn_module_defined=1 */ ;
    input \notGate[215]_keep ;
    output \notGate[216] ;
    
    wire \notGate[215]_keep  /* synthesis alspreserve=1 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(25[15:22])
    
    LUT4 I1 (.A(\notGate[215]_keep ), .B(\notGate[215]_keep ), .C(\notGate[215]_keep ), 
         .D(\notGate[215]_keep ), .Z(\notGate[216] )) /* synthesis syn_instantiated=1, lut_function=((!D !C !B !A)+(!D !C !B A)+(!D !C B !A)+(!D !C B A)+(!D C !B !A)+(!D C !B A)+(!D C B !A)+(!D C B A)), LSE_LINE_FILE_ID=3, LSE_LCOL=13, LSE_RCOL=44, LSE_LLINE=32, LSE_RLINE=32 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(11[2:53])
    defparam I1.init = 16'b0000000011111111;
    
endmodule
//
// Verilog Description of module inverter_U870
//

module inverter_U870 (\notGate[214]_keep , \notGate[215] ) /* synthesis syn_module_defined=1 */ ;
    input \notGate[214]_keep ;
    output \notGate[215] ;
    
    wire \notGate[214]_keep  /* synthesis alspreserve=1 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(25[15:22])
    
    LUT4 I1 (.A(\notGate[214]_keep ), .B(\notGate[214]_keep ), .C(\notGate[214]_keep ), 
         .D(\notGate[214]_keep ), .Z(\notGate[215] )) /* synthesis syn_instantiated=1, lut_function=((!D !C !B !A)+(!D !C !B A)+(!D !C B !A)+(!D !C B A)+(!D C !B !A)+(!D C !B A)+(!D C B !A)+(!D C B A)), LSE_LINE_FILE_ID=3, LSE_LCOL=13, LSE_RCOL=44, LSE_LLINE=32, LSE_RLINE=32 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(11[2:53])
    defparam I1.init = 16'b0000000011111111;
    
endmodule
//
// Verilog Description of module inverter_U871
//

module inverter_U871 (\notGate[213]_keep , \notGate[214] ) /* synthesis syn_module_defined=1 */ ;
    input \notGate[213]_keep ;
    output \notGate[214] ;
    
    wire \notGate[213]_keep  /* synthesis alspreserve=1 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(25[15:22])
    
    LUT4 I1 (.A(\notGate[213]_keep ), .B(\notGate[213]_keep ), .C(\notGate[213]_keep ), 
         .D(\notGate[213]_keep ), .Z(\notGate[214] )) /* synthesis syn_instantiated=1, lut_function=((!D !C !B !A)+(!D !C !B A)+(!D !C B !A)+(!D !C B A)+(!D C !B !A)+(!D C !B A)+(!D C B !A)+(!D C B A)), LSE_LINE_FILE_ID=3, LSE_LCOL=13, LSE_RCOL=44, LSE_LLINE=32, LSE_RLINE=32 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(11[2:53])
    defparam I1.init = 16'b0000000011111111;
    
endmodule
//
// Verilog Description of module inverter_U872
//

module inverter_U872 (\notGate[212]_keep , \notGate[213] ) /* synthesis syn_module_defined=1 */ ;
    input \notGate[212]_keep ;
    output \notGate[213] ;
    
    wire \notGate[212]_keep  /* synthesis alspreserve=1 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(25[15:22])
    
    LUT4 I1 (.A(\notGate[212]_keep ), .B(\notGate[212]_keep ), .C(\notGate[212]_keep ), 
         .D(\notGate[212]_keep ), .Z(\notGate[213] )) /* synthesis syn_instantiated=1, lut_function=((!D !C !B !A)+(!D !C !B A)+(!D !C B !A)+(!D !C B A)+(!D C !B !A)+(!D C !B A)+(!D C B !A)+(!D C B A)), LSE_LINE_FILE_ID=3, LSE_LCOL=13, LSE_RCOL=44, LSE_LLINE=32, LSE_RLINE=32 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(11[2:53])
    defparam I1.init = 16'b0000000011111111;
    
endmodule
//
// Verilog Description of module inverter_U873
//

module inverter_U873 (\notGate[211]_keep , \notGate[212] ) /* synthesis syn_module_defined=1 */ ;
    input \notGate[211]_keep ;
    output \notGate[212] ;
    
    wire \notGate[211]_keep  /* synthesis alspreserve=1 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(25[15:22])
    
    LUT4 I1 (.A(\notGate[211]_keep ), .B(\notGate[211]_keep ), .C(\notGate[211]_keep ), 
         .D(\notGate[211]_keep ), .Z(\notGate[212] )) /* synthesis syn_instantiated=1, lut_function=((!D !C !B !A)+(!D !C !B A)+(!D !C B !A)+(!D !C B A)+(!D C !B !A)+(!D C !B A)+(!D C B !A)+(!D C B A)), LSE_LINE_FILE_ID=3, LSE_LCOL=13, LSE_RCOL=44, LSE_LLINE=32, LSE_RLINE=32 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(11[2:53])
    defparam I1.init = 16'b0000000011111111;
    
endmodule
//
// Verilog Description of module inverter_U874
//

module inverter_U874 (\notGate[210]_keep , \notGate[211] ) /* synthesis syn_module_defined=1 */ ;
    input \notGate[210]_keep ;
    output \notGate[211] ;
    
    wire \notGate[210]_keep  /* synthesis alspreserve=1 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(25[15:22])
    
    LUT4 I1 (.A(\notGate[210]_keep ), .B(\notGate[210]_keep ), .C(\notGate[210]_keep ), 
         .D(\notGate[210]_keep ), .Z(\notGate[211] )) /* synthesis syn_instantiated=1, lut_function=((!D !C !B !A)+(!D !C !B A)+(!D !C B !A)+(!D !C B A)+(!D C !B !A)+(!D C !B A)+(!D C B !A)+(!D C B A)), LSE_LINE_FILE_ID=3, LSE_LCOL=13, LSE_RCOL=44, LSE_LLINE=32, LSE_RLINE=32 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(11[2:53])
    defparam I1.init = 16'b0000000011111111;
    
endmodule
//
// Verilog Description of module inverter_U875
//

module inverter_U875 (\notGate[209]_keep , \notGate[210] ) /* synthesis syn_module_defined=1 */ ;
    input \notGate[209]_keep ;
    output \notGate[210] ;
    
    wire \notGate[209]_keep  /* synthesis alspreserve=1 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(25[15:22])
    
    LUT4 I1 (.A(\notGate[209]_keep ), .B(\notGate[209]_keep ), .C(\notGate[209]_keep ), 
         .D(\notGate[209]_keep ), .Z(\notGate[210] )) /* synthesis syn_instantiated=1, lut_function=((!D !C !B !A)+(!D !C !B A)+(!D !C B !A)+(!D !C B A)+(!D C !B !A)+(!D C !B A)+(!D C B !A)+(!D C B A)), LSE_LINE_FILE_ID=3, LSE_LCOL=13, LSE_RCOL=44, LSE_LLINE=32, LSE_RLINE=32 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(11[2:53])
    defparam I1.init = 16'b0000000011111111;
    
endmodule
//
// Verilog Description of module inverter_U876
//

module inverter_U876 (\notGate[19]_keep , \notGate[20] ) /* synthesis syn_module_defined=1 */ ;
    input \notGate[19]_keep ;
    output \notGate[20] ;
    
    wire \notGate[19]_keep  /* synthesis alspreserve=1 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(25[15:22])
    
    LUT4 I1 (.A(\notGate[19]_keep ), .B(\notGate[19]_keep ), .C(\notGate[19]_keep ), 
         .D(\notGate[19]_keep ), .Z(\notGate[20] )) /* synthesis syn_instantiated=1, lut_function=((!D !C !B !A)+(!D !C !B A)+(!D !C B !A)+(!D !C B A)+(!D C !B !A)+(!D C !B A)+(!D C B !A)+(!D C B A)), LSE_LINE_FILE_ID=3, LSE_LCOL=13, LSE_RCOL=44, LSE_LLINE=32, LSE_RLINE=32 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(11[2:53])
    defparam I1.init = 16'b0000000011111111;
    
endmodule
//
// Verilog Description of module inverter_U877
//

module inverter_U877 (\notGate[208]_keep , \notGate[209] ) /* synthesis syn_module_defined=1 */ ;
    input \notGate[208]_keep ;
    output \notGate[209] ;
    
    wire \notGate[208]_keep  /* synthesis alspreserve=1 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(25[15:22])
    
    LUT4 I1 (.A(\notGate[208]_keep ), .B(\notGate[208]_keep ), .C(\notGate[208]_keep ), 
         .D(\notGate[208]_keep ), .Z(\notGate[209] )) /* synthesis syn_instantiated=1, lut_function=((!D !C !B !A)+(!D !C !B A)+(!D !C B !A)+(!D !C B A)+(!D C !B !A)+(!D C !B A)+(!D C B !A)+(!D C B A)), LSE_LINE_FILE_ID=3, LSE_LCOL=13, LSE_RCOL=44, LSE_LLINE=32, LSE_RLINE=32 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(11[2:53])
    defparam I1.init = 16'b0000000011111111;
    
endmodule
//
// Verilog Description of module inverter_U878
//

module inverter_U878 (\notGate[207]_keep , \notGate[208] ) /* synthesis syn_module_defined=1 */ ;
    input \notGate[207]_keep ;
    output \notGate[208] ;
    
    wire \notGate[207]_keep  /* synthesis alspreserve=1 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(25[15:22])
    
    LUT4 I1 (.A(\notGate[207]_keep ), .B(\notGate[207]_keep ), .C(\notGate[207]_keep ), 
         .D(\notGate[207]_keep ), .Z(\notGate[208] )) /* synthesis syn_instantiated=1, lut_function=((!D !C !B !A)+(!D !C !B A)+(!D !C B !A)+(!D !C B A)+(!D C !B !A)+(!D C !B A)+(!D C B !A)+(!D C B A)), LSE_LINE_FILE_ID=3, LSE_LCOL=13, LSE_RCOL=44, LSE_LLINE=32, LSE_RLINE=32 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(11[2:53])
    defparam I1.init = 16'b0000000011111111;
    
endmodule
//
// Verilog Description of module inverter_U879
//

module inverter_U879 (\notGate[206]_keep , \notGate[207] ) /* synthesis syn_module_defined=1 */ ;
    input \notGate[206]_keep ;
    output \notGate[207] ;
    
    wire \notGate[206]_keep  /* synthesis alspreserve=1 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(25[15:22])
    
    LUT4 I1 (.A(\notGate[206]_keep ), .B(\notGate[206]_keep ), .C(\notGate[206]_keep ), 
         .D(\notGate[206]_keep ), .Z(\notGate[207] )) /* synthesis syn_instantiated=1, lut_function=((!D !C !B !A)+(!D !C !B A)+(!D !C B !A)+(!D !C B A)+(!D C !B !A)+(!D C !B A)+(!D C B !A)+(!D C B A)), LSE_LINE_FILE_ID=3, LSE_LCOL=13, LSE_RCOL=44, LSE_LLINE=32, LSE_RLINE=32 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(11[2:53])
    defparam I1.init = 16'b0000000011111111;
    
endmodule
//
// Verilog Description of module inverter_U880
//

module inverter_U880 (\notGate[205]_keep , \notGate[206] ) /* synthesis syn_module_defined=1 */ ;
    input \notGate[205]_keep ;
    output \notGate[206] ;
    
    wire \notGate[205]_keep  /* synthesis alspreserve=1 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(25[15:22])
    
    LUT4 I1 (.A(\notGate[205]_keep ), .B(\notGate[205]_keep ), .C(\notGate[205]_keep ), 
         .D(\notGate[205]_keep ), .Z(\notGate[206] )) /* synthesis syn_instantiated=1, lut_function=((!D !C !B !A)+(!D !C !B A)+(!D !C B !A)+(!D !C B A)+(!D C !B !A)+(!D C !B A)+(!D C B !A)+(!D C B A)), LSE_LINE_FILE_ID=3, LSE_LCOL=13, LSE_RCOL=44, LSE_LLINE=32, LSE_RLINE=32 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(11[2:53])
    defparam I1.init = 16'b0000000011111111;
    
endmodule
//
// Verilog Description of module inverter_U881
//

module inverter_U881 (\notGate[204]_keep , \notGate[205] ) /* synthesis syn_module_defined=1 */ ;
    input \notGate[204]_keep ;
    output \notGate[205] ;
    
    wire \notGate[204]_keep  /* synthesis alspreserve=1 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(25[15:22])
    
    LUT4 I1 (.A(\notGate[204]_keep ), .B(\notGate[204]_keep ), .C(\notGate[204]_keep ), 
         .D(\notGate[204]_keep ), .Z(\notGate[205] )) /* synthesis syn_instantiated=1, lut_function=((!D !C !B !A)+(!D !C !B A)+(!D !C B !A)+(!D !C B A)+(!D C !B !A)+(!D C !B A)+(!D C B !A)+(!D C B A)), LSE_LINE_FILE_ID=3, LSE_LCOL=13, LSE_RCOL=44, LSE_LLINE=32, LSE_RLINE=32 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(11[2:53])
    defparam I1.init = 16'b0000000011111111;
    
endmodule
//
// Verilog Description of module inverter_U882
//

module inverter_U882 (\notGate[203]_keep , \notGate[204] ) /* synthesis syn_module_defined=1 */ ;
    input \notGate[203]_keep ;
    output \notGate[204] ;
    
    wire \notGate[203]_keep  /* synthesis alspreserve=1 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(25[15:22])
    
    LUT4 I1 (.A(\notGate[203]_keep ), .B(\notGate[203]_keep ), .C(\notGate[203]_keep ), 
         .D(\notGate[203]_keep ), .Z(\notGate[204] )) /* synthesis syn_instantiated=1, lut_function=((!D !C !B !A)+(!D !C !B A)+(!D !C B !A)+(!D !C B A)+(!D C !B !A)+(!D C !B A)+(!D C B !A)+(!D C B A)), LSE_LINE_FILE_ID=3, LSE_LCOL=13, LSE_RCOL=44, LSE_LLINE=32, LSE_RLINE=32 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(11[2:53])
    defparam I1.init = 16'b0000000011111111;
    
endmodule
//
// Verilog Description of module inverter_U883
//

module inverter_U883 (\notGate[202]_keep , \notGate[203] ) /* synthesis syn_module_defined=1 */ ;
    input \notGate[202]_keep ;
    output \notGate[203] ;
    
    wire \notGate[202]_keep  /* synthesis alspreserve=1 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(25[15:22])
    
    LUT4 I1 (.A(\notGate[202]_keep ), .B(\notGate[202]_keep ), .C(\notGate[202]_keep ), 
         .D(\notGate[202]_keep ), .Z(\notGate[203] )) /* synthesis syn_instantiated=1, lut_function=((!D !C !B !A)+(!D !C !B A)+(!D !C B !A)+(!D !C B A)+(!D C !B !A)+(!D C !B A)+(!D C B !A)+(!D C B A)), LSE_LINE_FILE_ID=3, LSE_LCOL=13, LSE_RCOL=44, LSE_LLINE=32, LSE_RLINE=32 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(11[2:53])
    defparam I1.init = 16'b0000000011111111;
    
endmodule
//
// Verilog Description of module inverter_U884
//

module inverter_U884 (\notGate[201]_keep , \notGate[202] ) /* synthesis syn_module_defined=1 */ ;
    input \notGate[201]_keep ;
    output \notGate[202] ;
    
    wire \notGate[201]_keep  /* synthesis alspreserve=1 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(25[15:22])
    
    LUT4 I1 (.A(\notGate[201]_keep ), .B(\notGate[201]_keep ), .C(\notGate[201]_keep ), 
         .D(\notGate[201]_keep ), .Z(\notGate[202] )) /* synthesis syn_instantiated=1, lut_function=((!D !C !B !A)+(!D !C !B A)+(!D !C B !A)+(!D !C B A)+(!D C !B !A)+(!D C !B A)+(!D C B !A)+(!D C B A)), LSE_LINE_FILE_ID=3, LSE_LCOL=13, LSE_RCOL=44, LSE_LLINE=32, LSE_RLINE=32 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(11[2:53])
    defparam I1.init = 16'b0000000011111111;
    
endmodule
//
// Verilog Description of module inverter_U885
//

module inverter_U885 (\notGate[200]_keep , \notGate[201] ) /* synthesis syn_module_defined=1 */ ;
    input \notGate[200]_keep ;
    output \notGate[201] ;
    
    wire \notGate[200]_keep  /* synthesis alspreserve=1 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(25[15:22])
    
    LUT4 I1 (.A(\notGate[200]_keep ), .B(\notGate[200]_keep ), .C(\notGate[200]_keep ), 
         .D(\notGate[200]_keep ), .Z(\notGate[201] )) /* synthesis syn_instantiated=1, lut_function=((!D !C !B !A)+(!D !C !B A)+(!D !C B !A)+(!D !C B A)+(!D C !B !A)+(!D C !B A)+(!D C B !A)+(!D C B A)), LSE_LINE_FILE_ID=3, LSE_LCOL=13, LSE_RCOL=44, LSE_LLINE=32, LSE_RLINE=32 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(11[2:53])
    defparam I1.init = 16'b0000000011111111;
    
endmodule
//
// Verilog Description of module inverter_U886
//

module inverter_U886 (\notGate[199]_keep , \notGate[200] ) /* synthesis syn_module_defined=1 */ ;
    input \notGate[199]_keep ;
    output \notGate[200] ;
    
    wire \notGate[199]_keep  /* synthesis alspreserve=1 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(25[15:22])
    
    LUT4 I1 (.A(\notGate[199]_keep ), .B(\notGate[199]_keep ), .C(\notGate[199]_keep ), 
         .D(\notGate[199]_keep ), .Z(\notGate[200] )) /* synthesis syn_instantiated=1, lut_function=((!D !C !B !A)+(!D !C !B A)+(!D !C B !A)+(!D !C B A)+(!D C !B !A)+(!D C !B A)+(!D C B !A)+(!D C B A)), LSE_LINE_FILE_ID=3, LSE_LCOL=13, LSE_RCOL=44, LSE_LLINE=32, LSE_RLINE=32 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(11[2:53])
    defparam I1.init = 16'b0000000011111111;
    
endmodule
//
// Verilog Description of module inverter_U887
//

module inverter_U887 (\notGate[0]_keep , \notGate[1] ) /* synthesis syn_module_defined=1 */ ;
    input \notGate[0]_keep ;
    output \notGate[1] ;
    
    wire \notGate[0]_keep  /* synthesis alspreserve=1 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(25[15:22])
    
    LUT4 I1 (.A(\notGate[0]_keep ), .B(\notGate[0]_keep ), .C(\notGate[0]_keep ), 
         .D(\notGate[0]_keep ), .Z(\notGate[1] )) /* synthesis syn_instantiated=1, lut_function=((!D !C !B !A)+(!D !C !B A)+(!D !C B !A)+(!D !C B A)+(!D C !B !A)+(!D C !B A)+(!D C B !A)+(!D C B A)), LSE_LINE_FILE_ID=3, LSE_LCOL=13, LSE_RCOL=44, LSE_LLINE=32, LSE_RLINE=32 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(11[2:53])
    defparam I1.init = 16'b0000000011111111;
    
endmodule
//
// Verilog Description of module inverter_U888
//

module inverter_U888 (\notGate[18]_keep , \notGate[19] ) /* synthesis syn_module_defined=1 */ ;
    input \notGate[18]_keep ;
    output \notGate[19] ;
    
    wire \notGate[18]_keep  /* synthesis alspreserve=1 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(25[15:22])
    
    LUT4 I1 (.A(\notGate[18]_keep ), .B(\notGate[18]_keep ), .C(\notGate[18]_keep ), 
         .D(\notGate[18]_keep ), .Z(\notGate[19] )) /* synthesis syn_instantiated=1, lut_function=((!D !C !B !A)+(!D !C !B A)+(!D !C B !A)+(!D !C B A)+(!D C !B !A)+(!D C !B A)+(!D C B !A)+(!D C B A)), LSE_LINE_FILE_ID=3, LSE_LCOL=13, LSE_RCOL=44, LSE_LLINE=32, LSE_RLINE=32 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(11[2:53])
    defparam I1.init = 16'b0000000011111111;
    
endmodule
//
// Verilog Description of module inverter_U889
//

module inverter_U889 (\notGate[198]_keep , \notGate[199] ) /* synthesis syn_module_defined=1 */ ;
    input \notGate[198]_keep ;
    output \notGate[199] ;
    
    wire \notGate[198]_keep  /* synthesis alspreserve=1 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(25[15:22])
    
    LUT4 I1 (.A(\notGate[198]_keep ), .B(\notGate[198]_keep ), .C(\notGate[198]_keep ), 
         .D(\notGate[198]_keep ), .Z(\notGate[199] )) /* synthesis syn_instantiated=1, lut_function=((!D !C !B !A)+(!D !C !B A)+(!D !C B !A)+(!D !C B A)+(!D C !B !A)+(!D C !B A)+(!D C B !A)+(!D C B A)), LSE_LINE_FILE_ID=3, LSE_LCOL=13, LSE_RCOL=44, LSE_LLINE=32, LSE_RLINE=32 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(11[2:53])
    defparam I1.init = 16'b0000000011111111;
    
endmodule
//
// Verilog Description of module inverter_U890
//

module inverter_U890 (\notGate[197]_keep , \notGate[198] ) /* synthesis syn_module_defined=1 */ ;
    input \notGate[197]_keep ;
    output \notGate[198] ;
    
    wire \notGate[197]_keep  /* synthesis alspreserve=1 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(25[15:22])
    
    LUT4 I1 (.A(\notGate[197]_keep ), .B(\notGate[197]_keep ), .C(\notGate[197]_keep ), 
         .D(\notGate[197]_keep ), .Z(\notGate[198] )) /* synthesis syn_instantiated=1, lut_function=((!D !C !B !A)+(!D !C !B A)+(!D !C B !A)+(!D !C B A)+(!D C !B !A)+(!D C !B A)+(!D C B !A)+(!D C B A)), LSE_LINE_FILE_ID=3, LSE_LCOL=13, LSE_RCOL=44, LSE_LLINE=32, LSE_RLINE=32 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(11[2:53])
    defparam I1.init = 16'b0000000011111111;
    
endmodule
//
// Verilog Description of module inverter_U891
//

module inverter_U891 (\notGate[196]_keep , \notGate[197] ) /* synthesis syn_module_defined=1 */ ;
    input \notGate[196]_keep ;
    output \notGate[197] ;
    
    wire \notGate[196]_keep  /* synthesis alspreserve=1 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(25[15:22])
    
    LUT4 I1 (.A(\notGate[196]_keep ), .B(\notGate[196]_keep ), .C(\notGate[196]_keep ), 
         .D(\notGate[196]_keep ), .Z(\notGate[197] )) /* synthesis syn_instantiated=1, lut_function=((!D !C !B !A)+(!D !C !B A)+(!D !C B !A)+(!D !C B A)+(!D C !B !A)+(!D C !B A)+(!D C B !A)+(!D C B A)), LSE_LINE_FILE_ID=3, LSE_LCOL=13, LSE_RCOL=44, LSE_LLINE=32, LSE_RLINE=32 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(11[2:53])
    defparam I1.init = 16'b0000000011111111;
    
endmodule
//
// Verilog Description of module inverter_U892
//

module inverter_U892 (\notGate[195]_keep , \notGate[196] ) /* synthesis syn_module_defined=1 */ ;
    input \notGate[195]_keep ;
    output \notGate[196] ;
    
    wire \notGate[195]_keep  /* synthesis alspreserve=1 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(25[15:22])
    
    LUT4 I1 (.A(\notGate[195]_keep ), .B(\notGate[195]_keep ), .C(\notGate[195]_keep ), 
         .D(\notGate[195]_keep ), .Z(\notGate[196] )) /* synthesis syn_instantiated=1, lut_function=((!D !C !B !A)+(!D !C !B A)+(!D !C B !A)+(!D !C B A)+(!D C !B !A)+(!D C !B A)+(!D C B !A)+(!D C B A)), LSE_LINE_FILE_ID=3, LSE_LCOL=13, LSE_RCOL=44, LSE_LLINE=32, LSE_RLINE=32 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(11[2:53])
    defparam I1.init = 16'b0000000011111111;
    
endmodule
//
// Verilog Description of module inverter_U893
//

module inverter_U893 (\notGate[194]_keep , \notGate[195] ) /* synthesis syn_module_defined=1 */ ;
    input \notGate[194]_keep ;
    output \notGate[195] ;
    
    wire \notGate[194]_keep  /* synthesis alspreserve=1 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(25[15:22])
    
    LUT4 I1 (.A(\notGate[194]_keep ), .B(\notGate[194]_keep ), .C(\notGate[194]_keep ), 
         .D(\notGate[194]_keep ), .Z(\notGate[195] )) /* synthesis syn_instantiated=1, lut_function=((!D !C !B !A)+(!D !C !B A)+(!D !C B !A)+(!D !C B A)+(!D C !B !A)+(!D C !B A)+(!D C B !A)+(!D C B A)), LSE_LINE_FILE_ID=3, LSE_LCOL=13, LSE_RCOL=44, LSE_LLINE=32, LSE_RLINE=32 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(11[2:53])
    defparam I1.init = 16'b0000000011111111;
    
endmodule
//
// Verilog Description of module inverter_U894
//

module inverter_U894 (\notGate[193]_keep , \notGate[194] ) /* synthesis syn_module_defined=1 */ ;
    input \notGate[193]_keep ;
    output \notGate[194] ;
    
    wire \notGate[193]_keep  /* synthesis alspreserve=1 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(25[15:22])
    
    LUT4 I1 (.A(\notGate[193]_keep ), .B(\notGate[193]_keep ), .C(\notGate[193]_keep ), 
         .D(\notGate[193]_keep ), .Z(\notGate[194] )) /* synthesis syn_instantiated=1, lut_function=((!D !C !B !A)+(!D !C !B A)+(!D !C B !A)+(!D !C B A)+(!D C !B !A)+(!D C !B A)+(!D C B !A)+(!D C B A)), LSE_LINE_FILE_ID=3, LSE_LCOL=13, LSE_RCOL=44, LSE_LLINE=32, LSE_RLINE=32 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(11[2:53])
    defparam I1.init = 16'b0000000011111111;
    
endmodule
//
// Verilog Description of module inverter_U895
//

module inverter_U895 (\notGate[192]_keep , \notGate[193] ) /* synthesis syn_module_defined=1 */ ;
    input \notGate[192]_keep ;
    output \notGate[193] ;
    
    wire \notGate[192]_keep  /* synthesis alspreserve=1 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(25[15:22])
    
    LUT4 I1 (.A(\notGate[192]_keep ), .B(\notGate[192]_keep ), .C(\notGate[192]_keep ), 
         .D(\notGate[192]_keep ), .Z(\notGate[193] )) /* synthesis syn_instantiated=1, lut_function=((!D !C !B !A)+(!D !C !B A)+(!D !C B !A)+(!D !C B A)+(!D C !B !A)+(!D C !B A)+(!D C B !A)+(!D C B A)), LSE_LINE_FILE_ID=3, LSE_LCOL=13, LSE_RCOL=44, LSE_LLINE=32, LSE_RLINE=32 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(11[2:53])
    defparam I1.init = 16'b0000000011111111;
    
endmodule
//
// Verilog Description of module inverter_U896
//

module inverter_U896 (\notGate[191]_keep , \notGate[192] ) /* synthesis syn_module_defined=1 */ ;
    input \notGate[191]_keep ;
    output \notGate[192] ;
    
    wire \notGate[191]_keep  /* synthesis alspreserve=1 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(25[15:22])
    
    LUT4 I1 (.A(\notGate[191]_keep ), .B(\notGate[191]_keep ), .C(\notGate[191]_keep ), 
         .D(\notGate[191]_keep ), .Z(\notGate[192] )) /* synthesis syn_instantiated=1, lut_function=((!D !C !B !A)+(!D !C !B A)+(!D !C B !A)+(!D !C B A)+(!D C !B !A)+(!D C !B A)+(!D C B !A)+(!D C B A)), LSE_LINE_FILE_ID=3, LSE_LCOL=13, LSE_RCOL=44, LSE_LLINE=32, LSE_RLINE=32 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(11[2:53])
    defparam I1.init = 16'b0000000011111111;
    
endmodule
//
// Verilog Description of module inverter_U897
//

module inverter_U897 (\notGate[190]_keep , \notGate[191] ) /* synthesis syn_module_defined=1 */ ;
    input \notGate[190]_keep ;
    output \notGate[191] ;
    
    wire \notGate[190]_keep  /* synthesis alspreserve=1 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(25[15:22])
    
    LUT4 I1 (.A(\notGate[190]_keep ), .B(\notGate[190]_keep ), .C(\notGate[190]_keep ), 
         .D(\notGate[190]_keep ), .Z(\notGate[191] )) /* synthesis syn_instantiated=1, lut_function=((!D !C !B !A)+(!D !C !B A)+(!D !C B !A)+(!D !C B A)+(!D C !B !A)+(!D C !B A)+(!D C B !A)+(!D C B A)), LSE_LINE_FILE_ID=3, LSE_LCOL=13, LSE_RCOL=44, LSE_LLINE=32, LSE_RLINE=32 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(11[2:53])
    defparam I1.init = 16'b0000000011111111;
    
endmodule
//
// Verilog Description of module inverter_U898
//

module inverter_U898 (\notGate[189]_keep , \notGate[190] ) /* synthesis syn_module_defined=1 */ ;
    input \notGate[189]_keep ;
    output \notGate[190] ;
    
    wire \notGate[189]_keep  /* synthesis alspreserve=1 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(25[15:22])
    
    LUT4 I1 (.A(\notGate[189]_keep ), .B(\notGate[189]_keep ), .C(\notGate[189]_keep ), 
         .D(\notGate[189]_keep ), .Z(\notGate[190] )) /* synthesis syn_instantiated=1, lut_function=((!D !C !B !A)+(!D !C !B A)+(!D !C B !A)+(!D !C B A)+(!D C !B !A)+(!D C !B A)+(!D C B !A)+(!D C B A)), LSE_LINE_FILE_ID=3, LSE_LCOL=13, LSE_RCOL=44, LSE_LLINE=32, LSE_RLINE=32 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(11[2:53])
    defparam I1.init = 16'b0000000011111111;
    
endmodule
//
// Verilog Description of module inverter_U899
//

module inverter_U899 (\notGate[17]_keep , \notGate[18] ) /* synthesis syn_module_defined=1 */ ;
    input \notGate[17]_keep ;
    output \notGate[18] ;
    
    wire \notGate[17]_keep  /* synthesis alspreserve=1 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(25[15:22])
    
    LUT4 I1 (.A(\notGate[17]_keep ), .B(\notGate[17]_keep ), .C(\notGate[17]_keep ), 
         .D(\notGate[17]_keep ), .Z(\notGate[18] )) /* synthesis syn_instantiated=1, lut_function=((!D !C !B !A)+(!D !C !B A)+(!D !C B !A)+(!D !C B A)+(!D C !B !A)+(!D C !B A)+(!D C B !A)+(!D C B A)), LSE_LINE_FILE_ID=3, LSE_LCOL=13, LSE_RCOL=44, LSE_LLINE=32, LSE_RLINE=32 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(11[2:53])
    defparam I1.init = 16'b0000000011111111;
    
endmodule
//
// Verilog Description of module inverter_U900
//

module inverter_U900 (\notGate[188]_keep , \notGate[189] ) /* synthesis syn_module_defined=1 */ ;
    input \notGate[188]_keep ;
    output \notGate[189] ;
    
    wire \notGate[188]_keep  /* synthesis alspreserve=1 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(25[15:22])
    
    LUT4 I1 (.A(\notGate[188]_keep ), .B(\notGate[188]_keep ), .C(\notGate[188]_keep ), 
         .D(\notGate[188]_keep ), .Z(\notGate[189] )) /* synthesis syn_instantiated=1, lut_function=((!D !C !B !A)+(!D !C !B A)+(!D !C B !A)+(!D !C B A)+(!D C !B !A)+(!D C !B A)+(!D C B !A)+(!D C B A)), LSE_LINE_FILE_ID=3, LSE_LCOL=13, LSE_RCOL=44, LSE_LLINE=32, LSE_RLINE=32 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(11[2:53])
    defparam I1.init = 16'b0000000011111111;
    
endmodule
//
// Verilog Description of module inverter_U901
//

module inverter_U901 (\notGate[187]_keep , \notGate[188] ) /* synthesis syn_module_defined=1 */ ;
    input \notGate[187]_keep ;
    output \notGate[188] ;
    
    wire \notGate[187]_keep  /* synthesis alspreserve=1 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(25[15:22])
    
    LUT4 I1 (.A(\notGate[187]_keep ), .B(\notGate[187]_keep ), .C(\notGate[187]_keep ), 
         .D(\notGate[187]_keep ), .Z(\notGate[188] )) /* synthesis syn_instantiated=1, lut_function=((!D !C !B !A)+(!D !C !B A)+(!D !C B !A)+(!D !C B A)+(!D C !B !A)+(!D C !B A)+(!D C B !A)+(!D C B A)), LSE_LINE_FILE_ID=3, LSE_LCOL=13, LSE_RCOL=44, LSE_LLINE=32, LSE_RLINE=32 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(11[2:53])
    defparam I1.init = 16'b0000000011111111;
    
endmodule
//
// Verilog Description of module inverter_U902
//

module inverter_U902 (\notGate[186]_keep , \notGate[187] ) /* synthesis syn_module_defined=1 */ ;
    input \notGate[186]_keep ;
    output \notGate[187] ;
    
    wire \notGate[186]_keep  /* synthesis alspreserve=1 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(25[15:22])
    
    LUT4 I1 (.A(\notGate[186]_keep ), .B(\notGate[186]_keep ), .C(\notGate[186]_keep ), 
         .D(\notGate[186]_keep ), .Z(\notGate[187] )) /* synthesis syn_instantiated=1, lut_function=((!D !C !B !A)+(!D !C !B A)+(!D !C B !A)+(!D !C B A)+(!D C !B !A)+(!D C !B A)+(!D C B !A)+(!D C B A)), LSE_LINE_FILE_ID=3, LSE_LCOL=13, LSE_RCOL=44, LSE_LLINE=32, LSE_RLINE=32 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(11[2:53])
    defparam I1.init = 16'b0000000011111111;
    
endmodule
//
// Verilog Description of module inverter_U903
//

module inverter_U903 (\notGate[185]_keep , \notGate[186] ) /* synthesis syn_module_defined=1 */ ;
    input \notGate[185]_keep ;
    output \notGate[186] ;
    
    wire \notGate[185]_keep  /* synthesis alspreserve=1 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(25[15:22])
    
    LUT4 I1 (.A(\notGate[185]_keep ), .B(\notGate[185]_keep ), .C(\notGate[185]_keep ), 
         .D(\notGate[185]_keep ), .Z(\notGate[186] )) /* synthesis syn_instantiated=1, lut_function=((!D !C !B !A)+(!D !C !B A)+(!D !C B !A)+(!D !C B A)+(!D C !B !A)+(!D C !B A)+(!D C B !A)+(!D C B A)), LSE_LINE_FILE_ID=3, LSE_LCOL=13, LSE_RCOL=44, LSE_LLINE=32, LSE_RLINE=32 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(11[2:53])
    defparam I1.init = 16'b0000000011111111;
    
endmodule
//
// Verilog Description of module inverter_U904
//

module inverter_U904 (\notGate[184]_keep , \notGate[185] ) /* synthesis syn_module_defined=1 */ ;
    input \notGate[184]_keep ;
    output \notGate[185] ;
    
    wire \notGate[184]_keep  /* synthesis alspreserve=1 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(25[15:22])
    
    LUT4 I1 (.A(\notGate[184]_keep ), .B(\notGate[184]_keep ), .C(\notGate[184]_keep ), 
         .D(\notGate[184]_keep ), .Z(\notGate[185] )) /* synthesis syn_instantiated=1, lut_function=((!D !C !B !A)+(!D !C !B A)+(!D !C B !A)+(!D !C B A)+(!D C !B !A)+(!D C !B A)+(!D C B !A)+(!D C B A)), LSE_LINE_FILE_ID=3, LSE_LCOL=13, LSE_RCOL=44, LSE_LLINE=32, LSE_RLINE=32 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(11[2:53])
    defparam I1.init = 16'b0000000011111111;
    
endmodule
//
// Verilog Description of module inverter_U905
//

module inverter_U905 (\notGate[183]_keep , \notGate[184] ) /* synthesis syn_module_defined=1 */ ;
    input \notGate[183]_keep ;
    output \notGate[184] ;
    
    wire \notGate[183]_keep  /* synthesis alspreserve=1 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(25[15:22])
    
    LUT4 I1 (.A(\notGate[183]_keep ), .B(\notGate[183]_keep ), .C(\notGate[183]_keep ), 
         .D(\notGate[183]_keep ), .Z(\notGate[184] )) /* synthesis syn_instantiated=1, lut_function=((!D !C !B !A)+(!D !C !B A)+(!D !C B !A)+(!D !C B A)+(!D C !B !A)+(!D C !B A)+(!D C B !A)+(!D C B A)), LSE_LINE_FILE_ID=3, LSE_LCOL=13, LSE_RCOL=44, LSE_LLINE=32, LSE_RLINE=32 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(11[2:53])
    defparam I1.init = 16'b0000000011111111;
    
endmodule
//
// Verilog Description of module inverter_U906
//

module inverter_U906 (\notGate[182]_keep , \notGate[183] ) /* synthesis syn_module_defined=1 */ ;
    input \notGate[182]_keep ;
    output \notGate[183] ;
    
    wire \notGate[182]_keep  /* synthesis alspreserve=1 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(25[15:22])
    
    LUT4 I1 (.A(\notGate[182]_keep ), .B(\notGate[182]_keep ), .C(\notGate[182]_keep ), 
         .D(\notGate[182]_keep ), .Z(\notGate[183] )) /* synthesis syn_instantiated=1, lut_function=((!D !C !B !A)+(!D !C !B A)+(!D !C B !A)+(!D !C B A)+(!D C !B !A)+(!D C !B A)+(!D C B !A)+(!D C B A)), LSE_LINE_FILE_ID=3, LSE_LCOL=13, LSE_RCOL=44, LSE_LLINE=32, LSE_RLINE=32 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(11[2:53])
    defparam I1.init = 16'b0000000011111111;
    
endmodule
//
// Verilog Description of module inverter_U907
//

module inverter_U907 (\notGate[181]_keep , \notGate[182] ) /* synthesis syn_module_defined=1 */ ;
    input \notGate[181]_keep ;
    output \notGate[182] ;
    
    wire \notGate[181]_keep  /* synthesis alspreserve=1 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(25[15:22])
    
    LUT4 I1 (.A(\notGate[181]_keep ), .B(\notGate[181]_keep ), .C(\notGate[181]_keep ), 
         .D(\notGate[181]_keep ), .Z(\notGate[182] )) /* synthesis syn_instantiated=1, lut_function=((!D !C !B !A)+(!D !C !B A)+(!D !C B !A)+(!D !C B A)+(!D C !B !A)+(!D C !B A)+(!D C B !A)+(!D C B A)), LSE_LINE_FILE_ID=3, LSE_LCOL=13, LSE_RCOL=44, LSE_LLINE=32, LSE_RLINE=32 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(11[2:53])
    defparam I1.init = 16'b0000000011111111;
    
endmodule
//
// Verilog Description of module inverter_U908
//

module inverter_U908 (\notGate[180]_keep , \notGate[181] ) /* synthesis syn_module_defined=1 */ ;
    input \notGate[180]_keep ;
    output \notGate[181] ;
    
    wire \notGate[180]_keep  /* synthesis alspreserve=1 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(25[15:22])
    
    LUT4 I1 (.A(\notGate[180]_keep ), .B(\notGate[180]_keep ), .C(\notGate[180]_keep ), 
         .D(\notGate[180]_keep ), .Z(\notGate[181] )) /* synthesis syn_instantiated=1, lut_function=((!D !C !B !A)+(!D !C !B A)+(!D !C B !A)+(!D !C B A)+(!D C !B !A)+(!D C !B A)+(!D C B !A)+(!D C B A)), LSE_LINE_FILE_ID=3, LSE_LCOL=13, LSE_RCOL=44, LSE_LLINE=32, LSE_RLINE=32 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(11[2:53])
    defparam I1.init = 16'b0000000011111111;
    
endmodule
//
// Verilog Description of module inverter_U909
//

module inverter_U909 (\notGate[179]_keep , \notGate[180] ) /* synthesis syn_module_defined=1 */ ;
    input \notGate[179]_keep ;
    output \notGate[180] ;
    
    wire \notGate[179]_keep  /* synthesis alspreserve=1 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(25[15:22])
    
    LUT4 I1 (.A(\notGate[179]_keep ), .B(\notGate[179]_keep ), .C(\notGate[179]_keep ), 
         .D(\notGate[179]_keep ), .Z(\notGate[180] )) /* synthesis syn_instantiated=1, lut_function=((!D !C !B !A)+(!D !C !B A)+(!D !C B !A)+(!D !C B A)+(!D C !B !A)+(!D C !B A)+(!D C B !A)+(!D C B A)), LSE_LINE_FILE_ID=3, LSE_LCOL=13, LSE_RCOL=44, LSE_LLINE=32, LSE_RLINE=32 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(11[2:53])
    defparam I1.init = 16'b0000000011111111;
    
endmodule
//
// Verilog Description of module inverter_U910
//

module inverter_U910 (\notGate[16]_keep , \notGate[17] ) /* synthesis syn_module_defined=1 */ ;
    input \notGate[16]_keep ;
    output \notGate[17] ;
    
    wire \notGate[16]_keep  /* synthesis alspreserve=1 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(25[15:22])
    
    LUT4 I1 (.A(\notGate[16]_keep ), .B(\notGate[16]_keep ), .C(\notGate[16]_keep ), 
         .D(\notGate[16]_keep ), .Z(\notGate[17] )) /* synthesis syn_instantiated=1, lut_function=((!D !C !B !A)+(!D !C !B A)+(!D !C B !A)+(!D !C B A)+(!D C !B !A)+(!D C !B A)+(!D C B !A)+(!D C B A)), LSE_LINE_FILE_ID=3, LSE_LCOL=13, LSE_RCOL=44, LSE_LLINE=32, LSE_RLINE=32 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(11[2:53])
    defparam I1.init = 16'b0000000011111111;
    
endmodule
//
// Verilog Description of module inverter_U911
//

module inverter_U911 (\notGate[178]_keep , \notGate[179] ) /* synthesis syn_module_defined=1 */ ;
    input \notGate[178]_keep ;
    output \notGate[179] ;
    
    wire \notGate[178]_keep  /* synthesis alspreserve=1 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(25[15:22])
    
    LUT4 I1 (.A(\notGate[178]_keep ), .B(\notGate[178]_keep ), .C(\notGate[178]_keep ), 
         .D(\notGate[178]_keep ), .Z(\notGate[179] )) /* synthesis syn_instantiated=1, lut_function=((!D !C !B !A)+(!D !C !B A)+(!D !C B !A)+(!D !C B A)+(!D C !B !A)+(!D C !B A)+(!D C B !A)+(!D C B A)), LSE_LINE_FILE_ID=3, LSE_LCOL=13, LSE_RCOL=44, LSE_LLINE=32, LSE_RLINE=32 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(11[2:53])
    defparam I1.init = 16'b0000000011111111;
    
endmodule
//
// Verilog Description of module inverter_U912
//

module inverter_U912 (\notGate[177]_keep , \notGate[178] ) /* synthesis syn_module_defined=1 */ ;
    input \notGate[177]_keep ;
    output \notGate[178] ;
    
    wire \notGate[177]_keep  /* synthesis alspreserve=1 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(25[15:22])
    
    LUT4 I1 (.A(\notGate[177]_keep ), .B(\notGate[177]_keep ), .C(\notGate[177]_keep ), 
         .D(\notGate[177]_keep ), .Z(\notGate[178] )) /* synthesis syn_instantiated=1, lut_function=((!D !C !B !A)+(!D !C !B A)+(!D !C B !A)+(!D !C B A)+(!D C !B !A)+(!D C !B A)+(!D C B !A)+(!D C B A)), LSE_LINE_FILE_ID=3, LSE_LCOL=13, LSE_RCOL=44, LSE_LLINE=32, LSE_RLINE=32 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(11[2:53])
    defparam I1.init = 16'b0000000011111111;
    
endmodule
//
// Verilog Description of module inverter_U913
//

module inverter_U913 (\notGate[176]_keep , \notGate[177] ) /* synthesis syn_module_defined=1 */ ;
    input \notGate[176]_keep ;
    output \notGate[177] ;
    
    wire \notGate[176]_keep  /* synthesis alspreserve=1 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(25[15:22])
    
    LUT4 I1 (.A(\notGate[176]_keep ), .B(\notGate[176]_keep ), .C(\notGate[176]_keep ), 
         .D(\notGate[176]_keep ), .Z(\notGate[177] )) /* synthesis syn_instantiated=1, lut_function=((!D !C !B !A)+(!D !C !B A)+(!D !C B !A)+(!D !C B A)+(!D C !B !A)+(!D C !B A)+(!D C B !A)+(!D C B A)), LSE_LINE_FILE_ID=3, LSE_LCOL=13, LSE_RCOL=44, LSE_LLINE=32, LSE_RLINE=32 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(11[2:53])
    defparam I1.init = 16'b0000000011111111;
    
endmodule
//
// Verilog Description of module inverter_U914
//

module inverter_U914 (\notGate[175]_keep , \notGate[176] ) /* synthesis syn_module_defined=1 */ ;
    input \notGate[175]_keep ;
    output \notGate[176] ;
    
    wire \notGate[175]_keep  /* synthesis alspreserve=1 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(25[15:22])
    
    LUT4 I1 (.A(\notGate[175]_keep ), .B(\notGate[175]_keep ), .C(\notGate[175]_keep ), 
         .D(\notGate[175]_keep ), .Z(\notGate[176] )) /* synthesis syn_instantiated=1, lut_function=((!D !C !B !A)+(!D !C !B A)+(!D !C B !A)+(!D !C B A)+(!D C !B !A)+(!D C !B A)+(!D C B !A)+(!D C B A)), LSE_LINE_FILE_ID=3, LSE_LCOL=13, LSE_RCOL=44, LSE_LLINE=32, LSE_RLINE=32 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(11[2:53])
    defparam I1.init = 16'b0000000011111111;
    
endmodule
//
// Verilog Description of module inverter_U915
//

module inverter_U915 (\notGate[174]_keep , \notGate[175] ) /* synthesis syn_module_defined=1 */ ;
    input \notGate[174]_keep ;
    output \notGate[175] ;
    
    wire \notGate[174]_keep  /* synthesis alspreserve=1 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(25[15:22])
    
    LUT4 I1 (.A(\notGate[174]_keep ), .B(\notGate[174]_keep ), .C(\notGate[174]_keep ), 
         .D(\notGate[174]_keep ), .Z(\notGate[175] )) /* synthesis syn_instantiated=1, lut_function=((!D !C !B !A)+(!D !C !B A)+(!D !C B !A)+(!D !C B A)+(!D C !B !A)+(!D C !B A)+(!D C B !A)+(!D C B A)), LSE_LINE_FILE_ID=3, LSE_LCOL=13, LSE_RCOL=44, LSE_LLINE=32, LSE_RLINE=32 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(11[2:53])
    defparam I1.init = 16'b0000000011111111;
    
endmodule
//
// Verilog Description of module inverter_U916
//

module inverter_U916 (\notGate[173]_keep , \notGate[174] ) /* synthesis syn_module_defined=1 */ ;
    input \notGate[173]_keep ;
    output \notGate[174] ;
    
    wire \notGate[173]_keep  /* synthesis alspreserve=1 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(25[15:22])
    
    LUT4 I1 (.A(\notGate[173]_keep ), .B(\notGate[173]_keep ), .C(\notGate[173]_keep ), 
         .D(\notGate[173]_keep ), .Z(\notGate[174] )) /* synthesis syn_instantiated=1, lut_function=((!D !C !B !A)+(!D !C !B A)+(!D !C B !A)+(!D !C B A)+(!D C !B !A)+(!D C !B A)+(!D C B !A)+(!D C B A)), LSE_LINE_FILE_ID=3, LSE_LCOL=13, LSE_RCOL=44, LSE_LLINE=32, LSE_RLINE=32 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(11[2:53])
    defparam I1.init = 16'b0000000011111111;
    
endmodule
//
// Verilog Description of module inverter_U917
//

module inverter_U917 (\notGate[172]_keep , \notGate[173] ) /* synthesis syn_module_defined=1 */ ;
    input \notGate[172]_keep ;
    output \notGate[173] ;
    
    wire \notGate[172]_keep  /* synthesis alspreserve=1 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(25[15:22])
    
    LUT4 I1 (.A(\notGate[172]_keep ), .B(\notGate[172]_keep ), .C(\notGate[172]_keep ), 
         .D(\notGate[172]_keep ), .Z(\notGate[173] )) /* synthesis syn_instantiated=1, lut_function=((!D !C !B !A)+(!D !C !B A)+(!D !C B !A)+(!D !C B A)+(!D C !B !A)+(!D C !B A)+(!D C B !A)+(!D C B A)), LSE_LINE_FILE_ID=3, LSE_LCOL=13, LSE_RCOL=44, LSE_LLINE=32, LSE_RLINE=32 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(11[2:53])
    defparam I1.init = 16'b0000000011111111;
    
endmodule
//
// Verilog Description of module inverter_U918
//

module inverter_U918 (\notGate[171]_keep , \notGate[172] ) /* synthesis syn_module_defined=1 */ ;
    input \notGate[171]_keep ;
    output \notGate[172] ;
    
    wire \notGate[171]_keep  /* synthesis alspreserve=1 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(25[15:22])
    
    LUT4 I1 (.A(\notGate[171]_keep ), .B(\notGate[171]_keep ), .C(\notGate[171]_keep ), 
         .D(\notGate[171]_keep ), .Z(\notGate[172] )) /* synthesis syn_instantiated=1, lut_function=((!D !C !B !A)+(!D !C !B A)+(!D !C B !A)+(!D !C B A)+(!D C !B !A)+(!D C !B A)+(!D C B !A)+(!D C B A)), LSE_LINE_FILE_ID=3, LSE_LCOL=13, LSE_RCOL=44, LSE_LLINE=32, LSE_RLINE=32 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(11[2:53])
    defparam I1.init = 16'b0000000011111111;
    
endmodule
//
// Verilog Description of module inverter_U919
//

module inverter_U919 (\notGate[170]_keep , \notGate[171] ) /* synthesis syn_module_defined=1 */ ;
    input \notGate[170]_keep ;
    output \notGate[171] ;
    
    wire \notGate[170]_keep  /* synthesis alspreserve=1 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(25[15:22])
    
    LUT4 I1 (.A(\notGate[170]_keep ), .B(\notGate[170]_keep ), .C(\notGate[170]_keep ), 
         .D(\notGate[170]_keep ), .Z(\notGate[171] )) /* synthesis syn_instantiated=1, lut_function=((!D !C !B !A)+(!D !C !B A)+(!D !C B !A)+(!D !C B A)+(!D C !B !A)+(!D C !B A)+(!D C B !A)+(!D C B A)), LSE_LINE_FILE_ID=3, LSE_LCOL=13, LSE_RCOL=44, LSE_LLINE=32, LSE_RLINE=32 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(11[2:53])
    defparam I1.init = 16'b0000000011111111;
    
endmodule
//
// Verilog Description of module inverter_U920
//

module inverter_U920 (\notGate[169]_keep , \notGate[170] ) /* synthesis syn_module_defined=1 */ ;
    input \notGate[169]_keep ;
    output \notGate[170] ;
    
    wire \notGate[169]_keep  /* synthesis alspreserve=1 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(25[15:22])
    
    LUT4 I1 (.A(\notGate[169]_keep ), .B(\notGate[169]_keep ), .C(\notGate[169]_keep ), 
         .D(\notGate[169]_keep ), .Z(\notGate[170] )) /* synthesis syn_instantiated=1, lut_function=((!D !C !B !A)+(!D !C !B A)+(!D !C B !A)+(!D !C B A)+(!D C !B !A)+(!D C !B A)+(!D C B !A)+(!D C B A)), LSE_LINE_FILE_ID=3, LSE_LCOL=13, LSE_RCOL=44, LSE_LLINE=32, LSE_RLINE=32 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(11[2:53])
    defparam I1.init = 16'b0000000011111111;
    
endmodule
//
// Verilog Description of module inverter_U921
//

module inverter_U921 (\notGate[15]_keep , \notGate[16] ) /* synthesis syn_module_defined=1 */ ;
    input \notGate[15]_keep ;
    output \notGate[16] ;
    
    wire \notGate[15]_keep  /* synthesis alspreserve=1 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(25[15:22])
    
    LUT4 I1 (.A(\notGate[15]_keep ), .B(\notGate[15]_keep ), .C(\notGate[15]_keep ), 
         .D(\notGate[15]_keep ), .Z(\notGate[16] )) /* synthesis syn_instantiated=1, lut_function=((!D !C !B !A)+(!D !C !B A)+(!D !C B !A)+(!D !C B A)+(!D C !B !A)+(!D C !B A)+(!D C B !A)+(!D C B A)), LSE_LINE_FILE_ID=3, LSE_LCOL=13, LSE_RCOL=44, LSE_LLINE=32, LSE_RLINE=32 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(11[2:53])
    defparam I1.init = 16'b0000000011111111;
    
endmodule
//
// Verilog Description of module inverter_U922
//

module inverter_U922 (\notGate[168]_keep , \notGate[169] ) /* synthesis syn_module_defined=1 */ ;
    input \notGate[168]_keep ;
    output \notGate[169] ;
    
    wire \notGate[168]_keep  /* synthesis alspreserve=1 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(25[15:22])
    
    LUT4 I1 (.A(\notGate[168]_keep ), .B(\notGate[168]_keep ), .C(\notGate[168]_keep ), 
         .D(\notGate[168]_keep ), .Z(\notGate[169] )) /* synthesis syn_instantiated=1, lut_function=((!D !C !B !A)+(!D !C !B A)+(!D !C B !A)+(!D !C B A)+(!D C !B !A)+(!D C !B A)+(!D C B !A)+(!D C B A)), LSE_LINE_FILE_ID=3, LSE_LCOL=13, LSE_RCOL=44, LSE_LLINE=32, LSE_RLINE=32 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(11[2:53])
    defparam I1.init = 16'b0000000011111111;
    
endmodule
//
// Verilog Description of module inverter_U923
//

module inverter_U923 (\notGate[167]_keep , \notGate[168] ) /* synthesis syn_module_defined=1 */ ;
    input \notGate[167]_keep ;
    output \notGate[168] ;
    
    wire \notGate[167]_keep  /* synthesis alspreserve=1 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(25[15:22])
    
    LUT4 I1 (.A(\notGate[167]_keep ), .B(\notGate[167]_keep ), .C(\notGate[167]_keep ), 
         .D(\notGate[167]_keep ), .Z(\notGate[168] )) /* synthesis syn_instantiated=1, lut_function=((!D !C !B !A)+(!D !C !B A)+(!D !C B !A)+(!D !C B A)+(!D C !B !A)+(!D C !B A)+(!D C B !A)+(!D C B A)), LSE_LINE_FILE_ID=3, LSE_LCOL=13, LSE_RCOL=44, LSE_LLINE=32, LSE_RLINE=32 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(11[2:53])
    defparam I1.init = 16'b0000000011111111;
    
endmodule
//
// Verilog Description of module inverter_U924
//

module inverter_U924 (\notGate[166]_keep , \notGate[167] ) /* synthesis syn_module_defined=1 */ ;
    input \notGate[166]_keep ;
    output \notGate[167] ;
    
    wire \notGate[166]_keep  /* synthesis alspreserve=1 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(25[15:22])
    
    LUT4 I1 (.A(\notGate[166]_keep ), .B(\notGate[166]_keep ), .C(\notGate[166]_keep ), 
         .D(\notGate[166]_keep ), .Z(\notGate[167] )) /* synthesis syn_instantiated=1, lut_function=((!D !C !B !A)+(!D !C !B A)+(!D !C B !A)+(!D !C B A)+(!D C !B !A)+(!D C !B A)+(!D C B !A)+(!D C B A)), LSE_LINE_FILE_ID=3, LSE_LCOL=13, LSE_RCOL=44, LSE_LLINE=32, LSE_RLINE=32 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(11[2:53])
    defparam I1.init = 16'b0000000011111111;
    
endmodule
//
// Verilog Description of module inverter_U925
//

module inverter_U925 (\notGate[165]_keep , \notGate[166] ) /* synthesis syn_module_defined=1 */ ;
    input \notGate[165]_keep ;
    output \notGate[166] ;
    
    wire \notGate[165]_keep  /* synthesis alspreserve=1 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(25[15:22])
    
    LUT4 I1 (.A(\notGate[165]_keep ), .B(\notGate[165]_keep ), .C(\notGate[165]_keep ), 
         .D(\notGate[165]_keep ), .Z(\notGate[166] )) /* synthesis syn_instantiated=1, lut_function=((!D !C !B !A)+(!D !C !B A)+(!D !C B !A)+(!D !C B A)+(!D C !B !A)+(!D C !B A)+(!D C B !A)+(!D C B A)), LSE_LINE_FILE_ID=3, LSE_LCOL=13, LSE_RCOL=44, LSE_LLINE=32, LSE_RLINE=32 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(11[2:53])
    defparam I1.init = 16'b0000000011111111;
    
endmodule
//
// Verilog Description of module inverter_U926
//

module inverter_U926 (\notGate[164]_keep , \notGate[165] ) /* synthesis syn_module_defined=1 */ ;
    input \notGate[164]_keep ;
    output \notGate[165] ;
    
    wire \notGate[164]_keep  /* synthesis alspreserve=1 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(25[15:22])
    
    LUT4 I1 (.A(\notGate[164]_keep ), .B(\notGate[164]_keep ), .C(\notGate[164]_keep ), 
         .D(\notGate[164]_keep ), .Z(\notGate[165] )) /* synthesis syn_instantiated=1, lut_function=((!D !C !B !A)+(!D !C !B A)+(!D !C B !A)+(!D !C B A)+(!D C !B !A)+(!D C !B A)+(!D C B !A)+(!D C B A)), LSE_LINE_FILE_ID=3, LSE_LCOL=13, LSE_RCOL=44, LSE_LLINE=32, LSE_RLINE=32 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(11[2:53])
    defparam I1.init = 16'b0000000011111111;
    
endmodule
//
// Verilog Description of module inverter_U927
//

module inverter_U927 (\notGate[163]_keep , \notGate[164] ) /* synthesis syn_module_defined=1 */ ;
    input \notGate[163]_keep ;
    output \notGate[164] ;
    
    wire \notGate[163]_keep  /* synthesis alspreserve=1 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(25[15:22])
    
    LUT4 I1 (.A(\notGate[163]_keep ), .B(\notGate[163]_keep ), .C(\notGate[163]_keep ), 
         .D(\notGate[163]_keep ), .Z(\notGate[164] )) /* synthesis syn_instantiated=1, lut_function=((!D !C !B !A)+(!D !C !B A)+(!D !C B !A)+(!D !C B A)+(!D C !B !A)+(!D C !B A)+(!D C B !A)+(!D C B A)), LSE_LINE_FILE_ID=3, LSE_LCOL=13, LSE_RCOL=44, LSE_LLINE=32, LSE_RLINE=32 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(11[2:53])
    defparam I1.init = 16'b0000000011111111;
    
endmodule
//
// Verilog Description of module inverter_U928
//

module inverter_U928 (\notGate[162]_keep , \notGate[163] ) /* synthesis syn_module_defined=1 */ ;
    input \notGate[162]_keep ;
    output \notGate[163] ;
    
    wire \notGate[162]_keep  /* synthesis alspreserve=1 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(25[15:22])
    
    LUT4 I1 (.A(\notGate[162]_keep ), .B(\notGate[162]_keep ), .C(\notGate[162]_keep ), 
         .D(\notGate[162]_keep ), .Z(\notGate[163] )) /* synthesis syn_instantiated=1, lut_function=((!D !C !B !A)+(!D !C !B A)+(!D !C B !A)+(!D !C B A)+(!D C !B !A)+(!D C !B A)+(!D C B !A)+(!D C B A)), LSE_LINE_FILE_ID=3, LSE_LCOL=13, LSE_RCOL=44, LSE_LLINE=32, LSE_RLINE=32 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(11[2:53])
    defparam I1.init = 16'b0000000011111111;
    
endmodule
//
// Verilog Description of module inverter_U929
//

module inverter_U929 (\notGate[161]_keep , \notGate[162] ) /* synthesis syn_module_defined=1 */ ;
    input \notGate[161]_keep ;
    output \notGate[162] ;
    
    wire \notGate[161]_keep  /* synthesis alspreserve=1 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(25[15:22])
    
    LUT4 I1 (.A(\notGate[161]_keep ), .B(\notGate[161]_keep ), .C(\notGate[161]_keep ), 
         .D(\notGate[161]_keep ), .Z(\notGate[162] )) /* synthesis syn_instantiated=1, lut_function=((!D !C !B !A)+(!D !C !B A)+(!D !C B !A)+(!D !C B A)+(!D C !B !A)+(!D C !B A)+(!D C B !A)+(!D C B A)), LSE_LINE_FILE_ID=3, LSE_LCOL=13, LSE_RCOL=44, LSE_LLINE=32, LSE_RLINE=32 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(11[2:53])
    defparam I1.init = 16'b0000000011111111;
    
endmodule
//
// Verilog Description of module inverter_U930
//

module inverter_U930 (\notGate[160]_keep , \notGate[161] ) /* synthesis syn_module_defined=1 */ ;
    input \notGate[160]_keep ;
    output \notGate[161] ;
    
    wire \notGate[160]_keep  /* synthesis alspreserve=1 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(25[15:22])
    
    LUT4 I1 (.A(\notGate[160]_keep ), .B(\notGate[160]_keep ), .C(\notGate[160]_keep ), 
         .D(\notGate[160]_keep ), .Z(\notGate[161] )) /* synthesis syn_instantiated=1, lut_function=((!D !C !B !A)+(!D !C !B A)+(!D !C B !A)+(!D !C B A)+(!D C !B !A)+(!D C !B A)+(!D C B !A)+(!D C B A)), LSE_LINE_FILE_ID=3, LSE_LCOL=13, LSE_RCOL=44, LSE_LLINE=32, LSE_RLINE=32 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(11[2:53])
    defparam I1.init = 16'b0000000011111111;
    
endmodule
//
// Verilog Description of module inverter_U931
//

module inverter_U931 (\notGate[159]_keep , \notGate[160] ) /* synthesis syn_module_defined=1 */ ;
    input \notGate[159]_keep ;
    output \notGate[160] ;
    
    wire \notGate[159]_keep  /* synthesis alspreserve=1 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(25[15:22])
    
    LUT4 I1 (.A(\notGate[159]_keep ), .B(\notGate[159]_keep ), .C(\notGate[159]_keep ), 
         .D(\notGate[159]_keep ), .Z(\notGate[160] )) /* synthesis syn_instantiated=1, lut_function=((!D !C !B !A)+(!D !C !B A)+(!D !C B !A)+(!D !C B A)+(!D C !B !A)+(!D C !B A)+(!D C B !A)+(!D C B A)), LSE_LINE_FILE_ID=3, LSE_LCOL=13, LSE_RCOL=44, LSE_LLINE=32, LSE_RLINE=32 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(11[2:53])
    defparam I1.init = 16'b0000000011111111;
    
endmodule
//
// Verilog Description of module inverter_U932
//

module inverter_U932 (\notGate[14]_keep , \notGate[15] ) /* synthesis syn_module_defined=1 */ ;
    input \notGate[14]_keep ;
    output \notGate[15] ;
    
    wire \notGate[14]_keep  /* synthesis alspreserve=1 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(25[15:22])
    
    LUT4 I1 (.A(\notGate[14]_keep ), .B(\notGate[14]_keep ), .C(\notGate[14]_keep ), 
         .D(\notGate[14]_keep ), .Z(\notGate[15] )) /* synthesis syn_instantiated=1, lut_function=((!D !C !B !A)+(!D !C !B A)+(!D !C B !A)+(!D !C B A)+(!D C !B !A)+(!D C !B A)+(!D C B !A)+(!D C B A)), LSE_LINE_FILE_ID=3, LSE_LCOL=13, LSE_RCOL=44, LSE_LLINE=32, LSE_RLINE=32 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(11[2:53])
    defparam I1.init = 16'b0000000011111111;
    
endmodule
//
// Verilog Description of module inverter_U933
//

module inverter_U933 (\notGate[158]_keep , \notGate[159] ) /* synthesis syn_module_defined=1 */ ;
    input \notGate[158]_keep ;
    output \notGate[159] ;
    
    wire \notGate[158]_keep  /* synthesis alspreserve=1 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(25[15:22])
    
    LUT4 I1 (.A(\notGate[158]_keep ), .B(\notGate[158]_keep ), .C(\notGate[158]_keep ), 
         .D(\notGate[158]_keep ), .Z(\notGate[159] )) /* synthesis syn_instantiated=1, lut_function=((!D !C !B !A)+(!D !C !B A)+(!D !C B !A)+(!D !C B A)+(!D C !B !A)+(!D C !B A)+(!D C B !A)+(!D C B A)), LSE_LINE_FILE_ID=3, LSE_LCOL=13, LSE_RCOL=44, LSE_LLINE=32, LSE_RLINE=32 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(11[2:53])
    defparam I1.init = 16'b0000000011111111;
    
endmodule
//
// Verilog Description of module inverter_U934
//

module inverter_U934 (\notGate[157]_keep , \notGate[158] ) /* synthesis syn_module_defined=1 */ ;
    input \notGate[157]_keep ;
    output \notGate[158] ;
    
    wire \notGate[157]_keep  /* synthesis alspreserve=1 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(25[15:22])
    
    LUT4 I1 (.A(\notGate[157]_keep ), .B(\notGate[157]_keep ), .C(\notGate[157]_keep ), 
         .D(\notGate[157]_keep ), .Z(\notGate[158] )) /* synthesis syn_instantiated=1, lut_function=((!D !C !B !A)+(!D !C !B A)+(!D !C B !A)+(!D !C B A)+(!D C !B !A)+(!D C !B A)+(!D C B !A)+(!D C B A)), LSE_LINE_FILE_ID=3, LSE_LCOL=13, LSE_RCOL=44, LSE_LLINE=32, LSE_RLINE=32 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(11[2:53])
    defparam I1.init = 16'b0000000011111111;
    
endmodule
//
// Verilog Description of module inverter_U935
//

module inverter_U935 (\notGate[156]_keep , \notGate[157] ) /* synthesis syn_module_defined=1 */ ;
    input \notGate[156]_keep ;
    output \notGate[157] ;
    
    wire \notGate[156]_keep  /* synthesis alspreserve=1 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(25[15:22])
    
    LUT4 I1 (.A(\notGate[156]_keep ), .B(\notGate[156]_keep ), .C(\notGate[156]_keep ), 
         .D(\notGate[156]_keep ), .Z(\notGate[157] )) /* synthesis syn_instantiated=1, lut_function=((!D !C !B !A)+(!D !C !B A)+(!D !C B !A)+(!D !C B A)+(!D C !B !A)+(!D C !B A)+(!D C B !A)+(!D C B A)), LSE_LINE_FILE_ID=3, LSE_LCOL=13, LSE_RCOL=44, LSE_LLINE=32, LSE_RLINE=32 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(11[2:53])
    defparam I1.init = 16'b0000000011111111;
    
endmodule
//
// Verilog Description of module inverter_U936
//

module inverter_U936 (\notGate[155]_keep , \notGate[156] ) /* synthesis syn_module_defined=1 */ ;
    input \notGate[155]_keep ;
    output \notGate[156] ;
    
    wire \notGate[155]_keep  /* synthesis alspreserve=1 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(25[15:22])
    
    LUT4 I1 (.A(\notGate[155]_keep ), .B(\notGate[155]_keep ), .C(\notGate[155]_keep ), 
         .D(\notGate[155]_keep ), .Z(\notGate[156] )) /* synthesis syn_instantiated=1, lut_function=((!D !C !B !A)+(!D !C !B A)+(!D !C B !A)+(!D !C B A)+(!D C !B !A)+(!D C !B A)+(!D C B !A)+(!D C B A)), LSE_LINE_FILE_ID=3, LSE_LCOL=13, LSE_RCOL=44, LSE_LLINE=32, LSE_RLINE=32 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(11[2:53])
    defparam I1.init = 16'b0000000011111111;
    
endmodule
//
// Verilog Description of module inverter_U937
//

module inverter_U937 (\notGate[154]_keep , \notGate[155] ) /* synthesis syn_module_defined=1 */ ;
    input \notGate[154]_keep ;
    output \notGate[155] ;
    
    wire \notGate[154]_keep  /* synthesis alspreserve=1 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(25[15:22])
    
    LUT4 I1 (.A(\notGate[154]_keep ), .B(\notGate[154]_keep ), .C(\notGate[154]_keep ), 
         .D(\notGate[154]_keep ), .Z(\notGate[155] )) /* synthesis syn_instantiated=1, lut_function=((!D !C !B !A)+(!D !C !B A)+(!D !C B !A)+(!D !C B A)+(!D C !B !A)+(!D C !B A)+(!D C B !A)+(!D C B A)), LSE_LINE_FILE_ID=3, LSE_LCOL=13, LSE_RCOL=44, LSE_LLINE=32, LSE_RLINE=32 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(11[2:53])
    defparam I1.init = 16'b0000000011111111;
    
endmodule
//
// Verilog Description of module inverter_U938
//

module inverter_U938 (\notGate[153]_keep , \notGate[154] ) /* synthesis syn_module_defined=1 */ ;
    input \notGate[153]_keep ;
    output \notGate[154] ;
    
    wire \notGate[153]_keep  /* synthesis alspreserve=1 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(25[15:22])
    
    LUT4 I1 (.A(\notGate[153]_keep ), .B(\notGate[153]_keep ), .C(\notGate[153]_keep ), 
         .D(\notGate[153]_keep ), .Z(\notGate[154] )) /* synthesis syn_instantiated=1, lut_function=((!D !C !B !A)+(!D !C !B A)+(!D !C B !A)+(!D !C B A)+(!D C !B !A)+(!D C !B A)+(!D C B !A)+(!D C B A)), LSE_LINE_FILE_ID=3, LSE_LCOL=13, LSE_RCOL=44, LSE_LLINE=32, LSE_RLINE=32 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(11[2:53])
    defparam I1.init = 16'b0000000011111111;
    
endmodule
//
// Verilog Description of module inverter_U939
//

module inverter_U939 (\notGate[152]_keep , \notGate[153] ) /* synthesis syn_module_defined=1 */ ;
    input \notGate[152]_keep ;
    output \notGate[153] ;
    
    wire \notGate[152]_keep  /* synthesis alspreserve=1 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(25[15:22])
    
    LUT4 I1 (.A(\notGate[152]_keep ), .B(\notGate[152]_keep ), .C(\notGate[152]_keep ), 
         .D(\notGate[152]_keep ), .Z(\notGate[153] )) /* synthesis syn_instantiated=1, lut_function=((!D !C !B !A)+(!D !C !B A)+(!D !C B !A)+(!D !C B A)+(!D C !B !A)+(!D C !B A)+(!D C B !A)+(!D C B A)), LSE_LINE_FILE_ID=3, LSE_LCOL=13, LSE_RCOL=44, LSE_LLINE=32, LSE_RLINE=32 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(11[2:53])
    defparam I1.init = 16'b0000000011111111;
    
endmodule
//
// Verilog Description of module inverter_U940
//

module inverter_U940 (\notGate[151]_keep , \notGate[152] ) /* synthesis syn_module_defined=1 */ ;
    input \notGate[151]_keep ;
    output \notGate[152] ;
    
    wire \notGate[151]_keep  /* synthesis alspreserve=1 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(25[15:22])
    
    LUT4 I1 (.A(\notGate[151]_keep ), .B(\notGate[151]_keep ), .C(\notGate[151]_keep ), 
         .D(\notGate[151]_keep ), .Z(\notGate[152] )) /* synthesis syn_instantiated=1, lut_function=((!D !C !B !A)+(!D !C !B A)+(!D !C B !A)+(!D !C B A)+(!D C !B !A)+(!D C !B A)+(!D C B !A)+(!D C B A)), LSE_LINE_FILE_ID=3, LSE_LCOL=13, LSE_RCOL=44, LSE_LLINE=32, LSE_RLINE=32 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(11[2:53])
    defparam I1.init = 16'b0000000011111111;
    
endmodule
//
// Verilog Description of module inverter_U941
//

module inverter_U941 (\notGate[150]_keep , \notGate[151] ) /* synthesis syn_module_defined=1 */ ;
    input \notGate[150]_keep ;
    output \notGate[151] ;
    
    wire \notGate[150]_keep  /* synthesis alspreserve=1 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(25[15:22])
    
    LUT4 I1 (.A(\notGate[150]_keep ), .B(\notGate[150]_keep ), .C(\notGate[150]_keep ), 
         .D(\notGate[150]_keep ), .Z(\notGate[151] )) /* synthesis syn_instantiated=1, lut_function=((!D !C !B !A)+(!D !C !B A)+(!D !C B !A)+(!D !C B A)+(!D C !B !A)+(!D C !B A)+(!D C B !A)+(!D C B A)), LSE_LINE_FILE_ID=3, LSE_LCOL=13, LSE_RCOL=44, LSE_LLINE=32, LSE_RLINE=32 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(11[2:53])
    defparam I1.init = 16'b0000000011111111;
    
endmodule
//
// Verilog Description of module inverter_U942
//

module inverter_U942 (\notGate[149]_keep , \notGate[150] ) /* synthesis syn_module_defined=1 */ ;
    input \notGate[149]_keep ;
    output \notGate[150] ;
    
    wire \notGate[149]_keep  /* synthesis alspreserve=1 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(25[15:22])
    
    LUT4 I1 (.A(\notGate[149]_keep ), .B(\notGate[149]_keep ), .C(\notGate[149]_keep ), 
         .D(\notGate[149]_keep ), .Z(\notGate[150] )) /* synthesis syn_instantiated=1, lut_function=((!D !C !B !A)+(!D !C !B A)+(!D !C B !A)+(!D !C B A)+(!D C !B !A)+(!D C !B A)+(!D C B !A)+(!D C B A)), LSE_LINE_FILE_ID=3, LSE_LCOL=13, LSE_RCOL=44, LSE_LLINE=32, LSE_RLINE=32 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(11[2:53])
    defparam I1.init = 16'b0000000011111111;
    
endmodule
//
// Verilog Description of module inverter_U943
//

module inverter_U943 (\notGate[13]_keep , \notGate[14] ) /* synthesis syn_module_defined=1 */ ;
    input \notGate[13]_keep ;
    output \notGate[14] ;
    
    wire \notGate[13]_keep  /* synthesis alspreserve=1 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(25[15:22])
    
    LUT4 I1 (.A(\notGate[13]_keep ), .B(\notGate[13]_keep ), .C(\notGate[13]_keep ), 
         .D(\notGate[13]_keep ), .Z(\notGate[14] )) /* synthesis syn_instantiated=1, lut_function=((!D !C !B !A)+(!D !C !B A)+(!D !C B !A)+(!D !C B A)+(!D C !B !A)+(!D C !B A)+(!D C B !A)+(!D C B A)), LSE_LINE_FILE_ID=3, LSE_LCOL=13, LSE_RCOL=44, LSE_LLINE=32, LSE_RLINE=32 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(11[2:53])
    defparam I1.init = 16'b0000000011111111;
    
endmodule
//
// Verilog Description of module inverter_U944
//

module inverter_U944 (\notGate[148]_keep , \notGate[149] ) /* synthesis syn_module_defined=1 */ ;
    input \notGate[148]_keep ;
    output \notGate[149] ;
    
    wire \notGate[148]_keep  /* synthesis alspreserve=1 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(25[15:22])
    
    LUT4 I1 (.A(\notGate[148]_keep ), .B(\notGate[148]_keep ), .C(\notGate[148]_keep ), 
         .D(\notGate[148]_keep ), .Z(\notGate[149] )) /* synthesis syn_instantiated=1, lut_function=((!D !C !B !A)+(!D !C !B A)+(!D !C B !A)+(!D !C B A)+(!D C !B !A)+(!D C !B A)+(!D C B !A)+(!D C B A)), LSE_LINE_FILE_ID=3, LSE_LCOL=13, LSE_RCOL=44, LSE_LLINE=32, LSE_RLINE=32 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(11[2:53])
    defparam I1.init = 16'b0000000011111111;
    
endmodule
//
// Verilog Description of module inverter_U945
//

module inverter_U945 (\notGate[147]_keep , \notGate[148] ) /* synthesis syn_module_defined=1 */ ;
    input \notGate[147]_keep ;
    output \notGate[148] ;
    
    wire \notGate[147]_keep  /* synthesis alspreserve=1 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(25[15:22])
    
    LUT4 I1 (.A(\notGate[147]_keep ), .B(\notGate[147]_keep ), .C(\notGate[147]_keep ), 
         .D(\notGate[147]_keep ), .Z(\notGate[148] )) /* synthesis syn_instantiated=1, lut_function=((!D !C !B !A)+(!D !C !B A)+(!D !C B !A)+(!D !C B A)+(!D C !B !A)+(!D C !B A)+(!D C B !A)+(!D C B A)), LSE_LINE_FILE_ID=3, LSE_LCOL=13, LSE_RCOL=44, LSE_LLINE=32, LSE_RLINE=32 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(11[2:53])
    defparam I1.init = 16'b0000000011111111;
    
endmodule
//
// Verilog Description of module inverter_U946
//

module inverter_U946 (\notGate[146]_keep , \notGate[147] ) /* synthesis syn_module_defined=1 */ ;
    input \notGate[146]_keep ;
    output \notGate[147] ;
    
    wire \notGate[146]_keep  /* synthesis alspreserve=1 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(25[15:22])
    
    LUT4 I1 (.A(\notGate[146]_keep ), .B(\notGate[146]_keep ), .C(\notGate[146]_keep ), 
         .D(\notGate[146]_keep ), .Z(\notGate[147] )) /* synthesis syn_instantiated=1, lut_function=((!D !C !B !A)+(!D !C !B A)+(!D !C B !A)+(!D !C B A)+(!D C !B !A)+(!D C !B A)+(!D C B !A)+(!D C B A)), LSE_LINE_FILE_ID=3, LSE_LCOL=13, LSE_RCOL=44, LSE_LLINE=32, LSE_RLINE=32 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(11[2:53])
    defparam I1.init = 16'b0000000011111111;
    
endmodule
//
// Verilog Description of module inverter_U947
//

module inverter_U947 (\notGate[145]_keep , \notGate[146] ) /* synthesis syn_module_defined=1 */ ;
    input \notGate[145]_keep ;
    output \notGate[146] ;
    
    wire \notGate[145]_keep  /* synthesis alspreserve=1 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(25[15:22])
    
    LUT4 I1 (.A(\notGate[145]_keep ), .B(\notGate[145]_keep ), .C(\notGate[145]_keep ), 
         .D(\notGate[145]_keep ), .Z(\notGate[146] )) /* synthesis syn_instantiated=1, lut_function=((!D !C !B !A)+(!D !C !B A)+(!D !C B !A)+(!D !C B A)+(!D C !B !A)+(!D C !B A)+(!D C B !A)+(!D C B A)), LSE_LINE_FILE_ID=3, LSE_LCOL=13, LSE_RCOL=44, LSE_LLINE=32, LSE_RLINE=32 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(11[2:53])
    defparam I1.init = 16'b0000000011111111;
    
endmodule
//
// Verilog Description of module inverter_U948
//

module inverter_U948 (\notGate[144]_keep , \notGate[145] ) /* synthesis syn_module_defined=1 */ ;
    input \notGate[144]_keep ;
    output \notGate[145] ;
    
    wire \notGate[144]_keep  /* synthesis alspreserve=1 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(25[15:22])
    
    LUT4 I1 (.A(\notGate[144]_keep ), .B(\notGate[144]_keep ), .C(\notGate[144]_keep ), 
         .D(\notGate[144]_keep ), .Z(\notGate[145] )) /* synthesis syn_instantiated=1, lut_function=((!D !C !B !A)+(!D !C !B A)+(!D !C B !A)+(!D !C B A)+(!D C !B !A)+(!D C !B A)+(!D C B !A)+(!D C B A)), LSE_LINE_FILE_ID=3, LSE_LCOL=13, LSE_RCOL=44, LSE_LLINE=32, LSE_RLINE=32 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(11[2:53])
    defparam I1.init = 16'b0000000011111111;
    
endmodule
//
// Verilog Description of module inverter_U949
//

module inverter_U949 (\notGate[143]_keep , \notGate[144] ) /* synthesis syn_module_defined=1 */ ;
    input \notGate[143]_keep ;
    output \notGate[144] ;
    
    wire \notGate[143]_keep  /* synthesis alspreserve=1 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(25[15:22])
    
    LUT4 I1 (.A(\notGate[143]_keep ), .B(\notGate[143]_keep ), .C(\notGate[143]_keep ), 
         .D(\notGate[143]_keep ), .Z(\notGate[144] )) /* synthesis syn_instantiated=1, lut_function=((!D !C !B !A)+(!D !C !B A)+(!D !C B !A)+(!D !C B A)+(!D C !B !A)+(!D C !B A)+(!D C B !A)+(!D C B A)), LSE_LINE_FILE_ID=3, LSE_LCOL=13, LSE_RCOL=44, LSE_LLINE=32, LSE_RLINE=32 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(11[2:53])
    defparam I1.init = 16'b0000000011111111;
    
endmodule
//
// Verilog Description of module inverter_U950
//

module inverter_U950 (\notGate[142]_keep , \notGate[143] ) /* synthesis syn_module_defined=1 */ ;
    input \notGate[142]_keep ;
    output \notGate[143] ;
    
    wire \notGate[142]_keep  /* synthesis alspreserve=1 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(25[15:22])
    
    LUT4 I1 (.A(\notGate[142]_keep ), .B(\notGate[142]_keep ), .C(\notGate[142]_keep ), 
         .D(\notGate[142]_keep ), .Z(\notGate[143] )) /* synthesis syn_instantiated=1, lut_function=((!D !C !B !A)+(!D !C !B A)+(!D !C B !A)+(!D !C B A)+(!D C !B !A)+(!D C !B A)+(!D C B !A)+(!D C B A)), LSE_LINE_FILE_ID=3, LSE_LCOL=13, LSE_RCOL=44, LSE_LLINE=32, LSE_RLINE=32 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(11[2:53])
    defparam I1.init = 16'b0000000011111111;
    
endmodule
//
// Verilog Description of module inverter_U951
//

module inverter_U951 (\notGate[141]_keep , \notGate[142] ) /* synthesis syn_module_defined=1 */ ;
    input \notGate[141]_keep ;
    output \notGate[142] ;
    
    wire \notGate[141]_keep  /* synthesis alspreserve=1 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(25[15:22])
    
    LUT4 I1 (.A(\notGate[141]_keep ), .B(\notGate[141]_keep ), .C(\notGate[141]_keep ), 
         .D(\notGate[141]_keep ), .Z(\notGate[142] )) /* synthesis syn_instantiated=1, lut_function=((!D !C !B !A)+(!D !C !B A)+(!D !C B !A)+(!D !C B A)+(!D C !B !A)+(!D C !B A)+(!D C B !A)+(!D C B A)), LSE_LINE_FILE_ID=3, LSE_LCOL=13, LSE_RCOL=44, LSE_LLINE=32, LSE_RLINE=32 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(11[2:53])
    defparam I1.init = 16'b0000000011111111;
    
endmodule
//
// Verilog Description of module inverter_U952
//

module inverter_U952 (\notGate[140]_keep , \notGate[141] ) /* synthesis syn_module_defined=1 */ ;
    input \notGate[140]_keep ;
    output \notGate[141] ;
    
    wire \notGate[140]_keep  /* synthesis alspreserve=1 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(25[15:22])
    
    LUT4 I1 (.A(\notGate[140]_keep ), .B(\notGate[140]_keep ), .C(\notGate[140]_keep ), 
         .D(\notGate[140]_keep ), .Z(\notGate[141] )) /* synthesis syn_instantiated=1, lut_function=((!D !C !B !A)+(!D !C !B A)+(!D !C B !A)+(!D !C B A)+(!D C !B !A)+(!D C !B A)+(!D C B !A)+(!D C B A)), LSE_LINE_FILE_ID=3, LSE_LCOL=13, LSE_RCOL=44, LSE_LLINE=32, LSE_RLINE=32 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(11[2:53])
    defparam I1.init = 16'b0000000011111111;
    
endmodule
//
// Verilog Description of module inverter_U953
//

module inverter_U953 (\notGate[139]_keep , \notGate[140] ) /* synthesis syn_module_defined=1 */ ;
    input \notGate[139]_keep ;
    output \notGate[140] ;
    
    wire \notGate[139]_keep  /* synthesis alspreserve=1 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(25[15:22])
    
    LUT4 I1 (.A(\notGate[139]_keep ), .B(\notGate[139]_keep ), .C(\notGate[139]_keep ), 
         .D(\notGate[139]_keep ), .Z(\notGate[140] )) /* synthesis syn_instantiated=1, lut_function=((!D !C !B !A)+(!D !C !B A)+(!D !C B !A)+(!D !C B A)+(!D C !B !A)+(!D C !B A)+(!D C B !A)+(!D C B A)), LSE_LINE_FILE_ID=3, LSE_LCOL=13, LSE_RCOL=44, LSE_LLINE=32, LSE_RLINE=32 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(11[2:53])
    defparam I1.init = 16'b0000000011111111;
    
endmodule
//
// Verilog Description of module inverter_U954
//

module inverter_U954 (\notGate[12]_keep , \notGate[13] ) /* synthesis syn_module_defined=1 */ ;
    input \notGate[12]_keep ;
    output \notGate[13] ;
    
    wire \notGate[12]_keep  /* synthesis alspreserve=1 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(25[15:22])
    
    LUT4 I1 (.A(\notGate[12]_keep ), .B(\notGate[12]_keep ), .C(\notGate[12]_keep ), 
         .D(\notGate[12]_keep ), .Z(\notGate[13] )) /* synthesis syn_instantiated=1, lut_function=((!D !C !B !A)+(!D !C !B A)+(!D !C B !A)+(!D !C B A)+(!D C !B !A)+(!D C !B A)+(!D C B !A)+(!D C B A)), LSE_LINE_FILE_ID=3, LSE_LCOL=13, LSE_RCOL=44, LSE_LLINE=32, LSE_RLINE=32 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(11[2:53])
    defparam I1.init = 16'b0000000011111111;
    
endmodule
//
// Verilog Description of module inverter_U955
//

module inverter_U955 (\notGate[138]_keep , \notGate[139] ) /* synthesis syn_module_defined=1 */ ;
    input \notGate[138]_keep ;
    output \notGate[139] ;
    
    wire \notGate[138]_keep  /* synthesis alspreserve=1 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(25[15:22])
    
    LUT4 I1 (.A(\notGate[138]_keep ), .B(\notGate[138]_keep ), .C(\notGate[138]_keep ), 
         .D(\notGate[138]_keep ), .Z(\notGate[139] )) /* synthesis syn_instantiated=1, lut_function=((!D !C !B !A)+(!D !C !B A)+(!D !C B !A)+(!D !C B A)+(!D C !B !A)+(!D C !B A)+(!D C B !A)+(!D C B A)), LSE_LINE_FILE_ID=3, LSE_LCOL=13, LSE_RCOL=44, LSE_LLINE=32, LSE_RLINE=32 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(11[2:53])
    defparam I1.init = 16'b0000000011111111;
    
endmodule
//
// Verilog Description of module inverter_U956
//

module inverter_U956 (\notGate[137]_keep , \notGate[138] ) /* synthesis syn_module_defined=1 */ ;
    input \notGate[137]_keep ;
    output \notGate[138] ;
    
    wire \notGate[137]_keep  /* synthesis alspreserve=1 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(25[15:22])
    
    LUT4 I1 (.A(\notGate[137]_keep ), .B(\notGate[137]_keep ), .C(\notGate[137]_keep ), 
         .D(\notGate[137]_keep ), .Z(\notGate[138] )) /* synthesis syn_instantiated=1, lut_function=((!D !C !B !A)+(!D !C !B A)+(!D !C B !A)+(!D !C B A)+(!D C !B !A)+(!D C !B A)+(!D C B !A)+(!D C B A)), LSE_LINE_FILE_ID=3, LSE_LCOL=13, LSE_RCOL=44, LSE_LLINE=32, LSE_RLINE=32 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(11[2:53])
    defparam I1.init = 16'b0000000011111111;
    
endmodule
//
// Verilog Description of module inverter_U957
//

module inverter_U957 (\notGate[136]_keep , \notGate[137] ) /* synthesis syn_module_defined=1 */ ;
    input \notGate[136]_keep ;
    output \notGate[137] ;
    
    wire \notGate[136]_keep  /* synthesis alspreserve=1 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(25[15:22])
    
    LUT4 I1 (.A(\notGate[136]_keep ), .B(\notGate[136]_keep ), .C(\notGate[136]_keep ), 
         .D(\notGate[136]_keep ), .Z(\notGate[137] )) /* synthesis syn_instantiated=1, lut_function=((!D !C !B !A)+(!D !C !B A)+(!D !C B !A)+(!D !C B A)+(!D C !B !A)+(!D C !B A)+(!D C B !A)+(!D C B A)), LSE_LINE_FILE_ID=3, LSE_LCOL=13, LSE_RCOL=44, LSE_LLINE=32, LSE_RLINE=32 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(11[2:53])
    defparam I1.init = 16'b0000000011111111;
    
endmodule
//
// Verilog Description of module inverter_U958
//

module inverter_U958 (\notGate[135]_keep , \notGate[136] ) /* synthesis syn_module_defined=1 */ ;
    input \notGate[135]_keep ;
    output \notGate[136] ;
    
    wire \notGate[135]_keep  /* synthesis alspreserve=1 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(25[15:22])
    
    LUT4 I1 (.A(\notGate[135]_keep ), .B(\notGate[135]_keep ), .C(\notGate[135]_keep ), 
         .D(\notGate[135]_keep ), .Z(\notGate[136] )) /* synthesis syn_instantiated=1, lut_function=((!D !C !B !A)+(!D !C !B A)+(!D !C B !A)+(!D !C B A)+(!D C !B !A)+(!D C !B A)+(!D C B !A)+(!D C B A)), LSE_LINE_FILE_ID=3, LSE_LCOL=13, LSE_RCOL=44, LSE_LLINE=32, LSE_RLINE=32 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(11[2:53])
    defparam I1.init = 16'b0000000011111111;
    
endmodule
//
// Verilog Description of module inverter_U959
//

module inverter_U959 (\notGate[134]_keep , \notGate[135] ) /* synthesis syn_module_defined=1 */ ;
    input \notGate[134]_keep ;
    output \notGate[135] ;
    
    wire \notGate[134]_keep  /* synthesis alspreserve=1 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(25[15:22])
    
    LUT4 I1 (.A(\notGate[134]_keep ), .B(\notGate[134]_keep ), .C(\notGate[134]_keep ), 
         .D(\notGate[134]_keep ), .Z(\notGate[135] )) /* synthesis syn_instantiated=1, lut_function=((!D !C !B !A)+(!D !C !B A)+(!D !C B !A)+(!D !C B A)+(!D C !B !A)+(!D C !B A)+(!D C B !A)+(!D C B A)), LSE_LINE_FILE_ID=3, LSE_LCOL=13, LSE_RCOL=44, LSE_LLINE=32, LSE_RLINE=32 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(11[2:53])
    defparam I1.init = 16'b0000000011111111;
    
endmodule
//
// Verilog Description of module inverter_U960
//

module inverter_U960 (\notGate[133]_keep , \notGate[134] ) /* synthesis syn_module_defined=1 */ ;
    input \notGate[133]_keep ;
    output \notGate[134] ;
    
    wire \notGate[133]_keep  /* synthesis alspreserve=1 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(25[15:22])
    
    LUT4 I1 (.A(\notGate[133]_keep ), .B(\notGate[133]_keep ), .C(\notGate[133]_keep ), 
         .D(\notGate[133]_keep ), .Z(\notGate[134] )) /* synthesis syn_instantiated=1, lut_function=((!D !C !B !A)+(!D !C !B A)+(!D !C B !A)+(!D !C B A)+(!D C !B !A)+(!D C !B A)+(!D C B !A)+(!D C B A)), LSE_LINE_FILE_ID=3, LSE_LCOL=13, LSE_RCOL=44, LSE_LLINE=32, LSE_RLINE=32 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(11[2:53])
    defparam I1.init = 16'b0000000011111111;
    
endmodule
//
// Verilog Description of module inverter_U961
//

module inverter_U961 (\notGate[132]_keep , \notGate[133] ) /* synthesis syn_module_defined=1 */ ;
    input \notGate[132]_keep ;
    output \notGate[133] ;
    
    wire \notGate[132]_keep  /* synthesis alspreserve=1 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(25[15:22])
    
    LUT4 I1 (.A(\notGate[132]_keep ), .B(\notGate[132]_keep ), .C(\notGate[132]_keep ), 
         .D(\notGate[132]_keep ), .Z(\notGate[133] )) /* synthesis syn_instantiated=1, lut_function=((!D !C !B !A)+(!D !C !B A)+(!D !C B !A)+(!D !C B A)+(!D C !B !A)+(!D C !B A)+(!D C B !A)+(!D C B A)), LSE_LINE_FILE_ID=3, LSE_LCOL=13, LSE_RCOL=44, LSE_LLINE=32, LSE_RLINE=32 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(11[2:53])
    defparam I1.init = 16'b0000000011111111;
    
endmodule
//
// Verilog Description of module inverter_U962
//

module inverter_U962 (\notGate[131]_keep , \notGate[132] ) /* synthesis syn_module_defined=1 */ ;
    input \notGate[131]_keep ;
    output \notGate[132] ;
    
    wire \notGate[131]_keep  /* synthesis alspreserve=1 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(25[15:22])
    
    LUT4 I1 (.A(\notGate[131]_keep ), .B(\notGate[131]_keep ), .C(\notGate[131]_keep ), 
         .D(\notGate[131]_keep ), .Z(\notGate[132] )) /* synthesis syn_instantiated=1, lut_function=((!D !C !B !A)+(!D !C !B A)+(!D !C B !A)+(!D !C B A)+(!D C !B !A)+(!D C !B A)+(!D C B !A)+(!D C B A)), LSE_LINE_FILE_ID=3, LSE_LCOL=13, LSE_RCOL=44, LSE_LLINE=32, LSE_RLINE=32 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(11[2:53])
    defparam I1.init = 16'b0000000011111111;
    
endmodule
//
// Verilog Description of module inverter_U963
//

module inverter_U963 (\notGate[130]_keep , \notGate[131] ) /* synthesis syn_module_defined=1 */ ;
    input \notGate[130]_keep ;
    output \notGate[131] ;
    
    wire \notGate[130]_keep  /* synthesis alspreserve=1 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(25[15:22])
    
    LUT4 I1 (.A(\notGate[130]_keep ), .B(\notGate[130]_keep ), .C(\notGate[130]_keep ), 
         .D(\notGate[130]_keep ), .Z(\notGate[131] )) /* synthesis syn_instantiated=1, lut_function=((!D !C !B !A)+(!D !C !B A)+(!D !C B !A)+(!D !C B A)+(!D C !B !A)+(!D C !B A)+(!D C B !A)+(!D C B A)), LSE_LINE_FILE_ID=3, LSE_LCOL=13, LSE_RCOL=44, LSE_LLINE=32, LSE_RLINE=32 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(11[2:53])
    defparam I1.init = 16'b0000000011111111;
    
endmodule
//
// Verilog Description of module inverter_U964
//

module inverter_U964 (\notGate[129]_keep , \notGate[130] ) /* synthesis syn_module_defined=1 */ ;
    input \notGate[129]_keep ;
    output \notGate[130] ;
    
    wire \notGate[129]_keep  /* synthesis alspreserve=1 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(25[15:22])
    
    LUT4 I1 (.A(\notGate[129]_keep ), .B(\notGate[129]_keep ), .C(\notGate[129]_keep ), 
         .D(\notGate[129]_keep ), .Z(\notGate[130] )) /* synthesis syn_instantiated=1, lut_function=((!D !C !B !A)+(!D !C !B A)+(!D !C B !A)+(!D !C B A)+(!D C !B !A)+(!D C !B A)+(!D C B !A)+(!D C B A)), LSE_LINE_FILE_ID=3, LSE_LCOL=13, LSE_RCOL=44, LSE_LLINE=32, LSE_RLINE=32 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(11[2:53])
    defparam I1.init = 16'b0000000011111111;
    
endmodule
//
// Verilog Description of module inverter_U965
//

module inverter_U965 (\notGate[11]_keep , \notGate[12] ) /* synthesis syn_module_defined=1 */ ;
    input \notGate[11]_keep ;
    output \notGate[12] ;
    
    wire \notGate[11]_keep  /* synthesis alspreserve=1 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(25[15:22])
    
    LUT4 I1 (.A(\notGate[11]_keep ), .B(\notGate[11]_keep ), .C(\notGate[11]_keep ), 
         .D(\notGate[11]_keep ), .Z(\notGate[12] )) /* synthesis syn_instantiated=1, lut_function=((!D !C !B !A)+(!D !C !B A)+(!D !C B !A)+(!D !C B A)+(!D C !B !A)+(!D C !B A)+(!D C B !A)+(!D C B A)), LSE_LINE_FILE_ID=3, LSE_LCOL=13, LSE_RCOL=44, LSE_LLINE=32, LSE_RLINE=32 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(11[2:53])
    defparam I1.init = 16'b0000000011111111;
    
endmodule
//
// Verilog Description of module inverter_U966
//

module inverter_U966 (\notGate[128]_keep , \notGate[129] ) /* synthesis syn_module_defined=1 */ ;
    input \notGate[128]_keep ;
    output \notGate[129] ;
    
    wire \notGate[128]_keep  /* synthesis alspreserve=1 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(25[15:22])
    
    LUT4 I1 (.A(\notGate[128]_keep ), .B(\notGate[128]_keep ), .C(\notGate[128]_keep ), 
         .D(\notGate[128]_keep ), .Z(\notGate[129] )) /* synthesis syn_instantiated=1, lut_function=((!D !C !B !A)+(!D !C !B A)+(!D !C B !A)+(!D !C B A)+(!D C !B !A)+(!D C !B A)+(!D C B !A)+(!D C B A)), LSE_LINE_FILE_ID=3, LSE_LCOL=13, LSE_RCOL=44, LSE_LLINE=32, LSE_RLINE=32 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(11[2:53])
    defparam I1.init = 16'b0000000011111111;
    
endmodule
//
// Verilog Description of module inverter_U967
//

module inverter_U967 (\notGate[127]_keep , \notGate[128] ) /* synthesis syn_module_defined=1 */ ;
    input \notGate[127]_keep ;
    output \notGate[128] ;
    
    wire \notGate[127]_keep  /* synthesis alspreserve=1 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(25[15:22])
    
    LUT4 I1 (.A(\notGate[127]_keep ), .B(\notGate[127]_keep ), .C(\notGate[127]_keep ), 
         .D(\notGate[127]_keep ), .Z(\notGate[128] )) /* synthesis syn_instantiated=1, lut_function=((!D !C !B !A)+(!D !C !B A)+(!D !C B !A)+(!D !C B A)+(!D C !B !A)+(!D C !B A)+(!D C B !A)+(!D C B A)), LSE_LINE_FILE_ID=3, LSE_LCOL=13, LSE_RCOL=44, LSE_LLINE=32, LSE_RLINE=32 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(11[2:53])
    defparam I1.init = 16'b0000000011111111;
    
endmodule
//
// Verilog Description of module inverter_U968
//

module inverter_U968 (\notGate[126]_keep , \notGate[127] ) /* synthesis syn_module_defined=1 */ ;
    input \notGate[126]_keep ;
    output \notGate[127] ;
    
    wire \notGate[126]_keep  /* synthesis alspreserve=1 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(25[15:22])
    
    LUT4 I1 (.A(\notGate[126]_keep ), .B(\notGate[126]_keep ), .C(\notGate[126]_keep ), 
         .D(\notGate[126]_keep ), .Z(\notGate[127] )) /* synthesis syn_instantiated=1, lut_function=((!D !C !B !A)+(!D !C !B A)+(!D !C B !A)+(!D !C B A)+(!D C !B !A)+(!D C !B A)+(!D C B !A)+(!D C B A)), LSE_LINE_FILE_ID=3, LSE_LCOL=13, LSE_RCOL=44, LSE_LLINE=32, LSE_RLINE=32 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(11[2:53])
    defparam I1.init = 16'b0000000011111111;
    
endmodule
//
// Verilog Description of module inverter_U969
//

module inverter_U969 (\notGate[125]_keep , \notGate[126] ) /* synthesis syn_module_defined=1 */ ;
    input \notGate[125]_keep ;
    output \notGate[126] ;
    
    wire \notGate[125]_keep  /* synthesis alspreserve=1 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(25[15:22])
    
    LUT4 I1 (.A(\notGate[125]_keep ), .B(\notGate[125]_keep ), .C(\notGate[125]_keep ), 
         .D(\notGate[125]_keep ), .Z(\notGate[126] )) /* synthesis syn_instantiated=1, lut_function=((!D !C !B !A)+(!D !C !B A)+(!D !C B !A)+(!D !C B A)+(!D C !B !A)+(!D C !B A)+(!D C B !A)+(!D C B A)), LSE_LINE_FILE_ID=3, LSE_LCOL=13, LSE_RCOL=44, LSE_LLINE=32, LSE_RLINE=32 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(11[2:53])
    defparam I1.init = 16'b0000000011111111;
    
endmodule
//
// Verilog Description of module inverter_U970
//

module inverter_U970 (\notGate[124]_keep , \notGate[125] ) /* synthesis syn_module_defined=1 */ ;
    input \notGate[124]_keep ;
    output \notGate[125] ;
    
    wire \notGate[124]_keep  /* synthesis alspreserve=1 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(25[15:22])
    
    LUT4 I1 (.A(\notGate[124]_keep ), .B(\notGate[124]_keep ), .C(\notGate[124]_keep ), 
         .D(\notGate[124]_keep ), .Z(\notGate[125] )) /* synthesis syn_instantiated=1, lut_function=((!D !C !B !A)+(!D !C !B A)+(!D !C B !A)+(!D !C B A)+(!D C !B !A)+(!D C !B A)+(!D C B !A)+(!D C B A)), LSE_LINE_FILE_ID=3, LSE_LCOL=13, LSE_RCOL=44, LSE_LLINE=32, LSE_RLINE=32 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(11[2:53])
    defparam I1.init = 16'b0000000011111111;
    
endmodule
//
// Verilog Description of module inverter_U971
//

module inverter_U971 (\notGate[123]_keep , \notGate[124] ) /* synthesis syn_module_defined=1 */ ;
    input \notGate[123]_keep ;
    output \notGate[124] ;
    
    wire \notGate[123]_keep  /* synthesis alspreserve=1 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(25[15:22])
    
    LUT4 I1 (.A(\notGate[123]_keep ), .B(\notGate[123]_keep ), .C(\notGate[123]_keep ), 
         .D(\notGate[123]_keep ), .Z(\notGate[124] )) /* synthesis syn_instantiated=1, lut_function=((!D !C !B !A)+(!D !C !B A)+(!D !C B !A)+(!D !C B A)+(!D C !B !A)+(!D C !B A)+(!D C B !A)+(!D C B A)), LSE_LINE_FILE_ID=3, LSE_LCOL=13, LSE_RCOL=44, LSE_LLINE=32, LSE_RLINE=32 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(11[2:53])
    defparam I1.init = 16'b0000000011111111;
    
endmodule
//
// Verilog Description of module inverter_U972
//

module inverter_U972 (\notGate[122]_keep , \notGate[123] ) /* synthesis syn_module_defined=1 */ ;
    input \notGate[122]_keep ;
    output \notGate[123] ;
    
    wire \notGate[122]_keep  /* synthesis alspreserve=1 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(25[15:22])
    
    LUT4 I1 (.A(\notGate[122]_keep ), .B(\notGate[122]_keep ), .C(\notGate[122]_keep ), 
         .D(\notGate[122]_keep ), .Z(\notGate[123] )) /* synthesis syn_instantiated=1, lut_function=((!D !C !B !A)+(!D !C !B A)+(!D !C B !A)+(!D !C B A)+(!D C !B !A)+(!D C !B A)+(!D C B !A)+(!D C B A)), LSE_LINE_FILE_ID=3, LSE_LCOL=13, LSE_RCOL=44, LSE_LLINE=32, LSE_RLINE=32 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(11[2:53])
    defparam I1.init = 16'b0000000011111111;
    
endmodule
//
// Verilog Description of module inverter_U973
//

module inverter_U973 (\notGate[121]_keep , \notGate[122] ) /* synthesis syn_module_defined=1 */ ;
    input \notGate[121]_keep ;
    output \notGate[122] ;
    
    wire \notGate[121]_keep  /* synthesis alspreserve=1 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(25[15:22])
    
    LUT4 I1 (.A(\notGate[121]_keep ), .B(\notGate[121]_keep ), .C(\notGate[121]_keep ), 
         .D(\notGate[121]_keep ), .Z(\notGate[122] )) /* synthesis syn_instantiated=1, lut_function=((!D !C !B !A)+(!D !C !B A)+(!D !C B !A)+(!D !C B A)+(!D C !B !A)+(!D C !B A)+(!D C B !A)+(!D C B A)), LSE_LINE_FILE_ID=3, LSE_LCOL=13, LSE_RCOL=44, LSE_LLINE=32, LSE_RLINE=32 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(11[2:53])
    defparam I1.init = 16'b0000000011111111;
    
endmodule
//
// Verilog Description of module inverter_U974
//

module inverter_U974 (\notGate[120]_keep , \notGate[121] ) /* synthesis syn_module_defined=1 */ ;
    input \notGate[120]_keep ;
    output \notGate[121] ;
    
    wire \notGate[120]_keep  /* synthesis alspreserve=1 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(25[15:22])
    
    LUT4 I1 (.A(\notGate[120]_keep ), .B(\notGate[120]_keep ), .C(\notGate[120]_keep ), 
         .D(\notGate[120]_keep ), .Z(\notGate[121] )) /* synthesis syn_instantiated=1, lut_function=((!D !C !B !A)+(!D !C !B A)+(!D !C B !A)+(!D !C B A)+(!D C !B !A)+(!D C !B A)+(!D C B !A)+(!D C B A)), LSE_LINE_FILE_ID=3, LSE_LCOL=13, LSE_RCOL=44, LSE_LLINE=32, LSE_RLINE=32 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(11[2:53])
    defparam I1.init = 16'b0000000011111111;
    
endmodule
//
// Verilog Description of module inverter_U975
//

module inverter_U975 (\notGate[119]_keep , \notGate[120] ) /* synthesis syn_module_defined=1 */ ;
    input \notGate[119]_keep ;
    output \notGate[120] ;
    
    wire \notGate[119]_keep  /* synthesis alspreserve=1 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(25[15:22])
    
    LUT4 I1 (.A(\notGate[119]_keep ), .B(\notGate[119]_keep ), .C(\notGate[119]_keep ), 
         .D(\notGate[119]_keep ), .Z(\notGate[120] )) /* synthesis syn_instantiated=1, lut_function=((!D !C !B !A)+(!D !C !B A)+(!D !C B !A)+(!D !C B A)+(!D C !B !A)+(!D C !B A)+(!D C B !A)+(!D C B A)), LSE_LINE_FILE_ID=3, LSE_LCOL=13, LSE_RCOL=44, LSE_LLINE=32, LSE_RLINE=32 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(11[2:53])
    defparam I1.init = 16'b0000000011111111;
    
endmodule
//
// Verilog Description of module inverter_U976
//

module inverter_U976 (\notGate[10]_keep , \notGate[11] ) /* synthesis syn_module_defined=1 */ ;
    input \notGate[10]_keep ;
    output \notGate[11] ;
    
    wire \notGate[10]_keep  /* synthesis alspreserve=1 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(25[15:22])
    
    LUT4 I1 (.A(\notGate[10]_keep ), .B(\notGate[10]_keep ), .C(\notGate[10]_keep ), 
         .D(\notGate[10]_keep ), .Z(\notGate[11] )) /* synthesis syn_instantiated=1, lut_function=((!D !C !B !A)+(!D !C !B A)+(!D !C B !A)+(!D !C B A)+(!D C !B !A)+(!D C !B A)+(!D C B !A)+(!D C B A)), LSE_LINE_FILE_ID=3, LSE_LCOL=13, LSE_RCOL=44, LSE_LLINE=32, LSE_RLINE=32 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(11[2:53])
    defparam I1.init = 16'b0000000011111111;
    
endmodule
//
// Verilog Description of module inverter_U977
//

module inverter_U977 (\notGate[118]_keep , \notGate[119] ) /* synthesis syn_module_defined=1 */ ;
    input \notGate[118]_keep ;
    output \notGate[119] ;
    
    wire \notGate[118]_keep  /* synthesis alspreserve=1 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(25[15:22])
    
    LUT4 I1 (.A(\notGate[118]_keep ), .B(\notGate[118]_keep ), .C(\notGate[118]_keep ), 
         .D(\notGate[118]_keep ), .Z(\notGate[119] )) /* synthesis syn_instantiated=1, lut_function=((!D !C !B !A)+(!D !C !B A)+(!D !C B !A)+(!D !C B A)+(!D C !B !A)+(!D C !B A)+(!D C B !A)+(!D C B A)), LSE_LINE_FILE_ID=3, LSE_LCOL=13, LSE_RCOL=44, LSE_LLINE=32, LSE_RLINE=32 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(11[2:53])
    defparam I1.init = 16'b0000000011111111;
    
endmodule
//
// Verilog Description of module inverter_U978
//

module inverter_U978 (\notGate[117]_keep , \notGate[118] ) /* synthesis syn_module_defined=1 */ ;
    input \notGate[117]_keep ;
    output \notGate[118] ;
    
    wire \notGate[117]_keep  /* synthesis alspreserve=1 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(25[15:22])
    
    LUT4 I1 (.A(\notGate[117]_keep ), .B(\notGate[117]_keep ), .C(\notGate[117]_keep ), 
         .D(\notGate[117]_keep ), .Z(\notGate[118] )) /* synthesis syn_instantiated=1, lut_function=((!D !C !B !A)+(!D !C !B A)+(!D !C B !A)+(!D !C B A)+(!D C !B !A)+(!D C !B A)+(!D C B !A)+(!D C B A)), LSE_LINE_FILE_ID=3, LSE_LCOL=13, LSE_RCOL=44, LSE_LLINE=32, LSE_RLINE=32 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(11[2:53])
    defparam I1.init = 16'b0000000011111111;
    
endmodule
//
// Verilog Description of module inverter_U979
//

module inverter_U979 (\notGate[116]_keep , \notGate[117] ) /* synthesis syn_module_defined=1 */ ;
    input \notGate[116]_keep ;
    output \notGate[117] ;
    
    wire \notGate[116]_keep  /* synthesis alspreserve=1 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(25[15:22])
    
    LUT4 I1 (.A(\notGate[116]_keep ), .B(\notGate[116]_keep ), .C(\notGate[116]_keep ), 
         .D(\notGate[116]_keep ), .Z(\notGate[117] )) /* synthesis syn_instantiated=1, lut_function=((!D !C !B !A)+(!D !C !B A)+(!D !C B !A)+(!D !C B A)+(!D C !B !A)+(!D C !B A)+(!D C B !A)+(!D C B A)), LSE_LINE_FILE_ID=3, LSE_LCOL=13, LSE_RCOL=44, LSE_LLINE=32, LSE_RLINE=32 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(11[2:53])
    defparam I1.init = 16'b0000000011111111;
    
endmodule
//
// Verilog Description of module inverter_U980
//

module inverter_U980 (\notGate[115]_keep , \notGate[116] ) /* synthesis syn_module_defined=1 */ ;
    input \notGate[115]_keep ;
    output \notGate[116] ;
    
    wire \notGate[115]_keep  /* synthesis alspreserve=1 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(25[15:22])
    
    LUT4 I1 (.A(\notGate[115]_keep ), .B(\notGate[115]_keep ), .C(\notGate[115]_keep ), 
         .D(\notGate[115]_keep ), .Z(\notGate[116] )) /* synthesis syn_instantiated=1, lut_function=((!D !C !B !A)+(!D !C !B A)+(!D !C B !A)+(!D !C B A)+(!D C !B !A)+(!D C !B A)+(!D C B !A)+(!D C B A)), LSE_LINE_FILE_ID=3, LSE_LCOL=13, LSE_RCOL=44, LSE_LLINE=32, LSE_RLINE=32 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(11[2:53])
    defparam I1.init = 16'b0000000011111111;
    
endmodule
//
// Verilog Description of module inverter_U981
//

module inverter_U981 (\notGate[114]_keep , \notGate[115] ) /* synthesis syn_module_defined=1 */ ;
    input \notGate[114]_keep ;
    output \notGate[115] ;
    
    wire \notGate[114]_keep  /* synthesis alspreserve=1 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(25[15:22])
    
    LUT4 I1 (.A(\notGate[114]_keep ), .B(\notGate[114]_keep ), .C(\notGate[114]_keep ), 
         .D(\notGate[114]_keep ), .Z(\notGate[115] )) /* synthesis syn_instantiated=1, lut_function=((!D !C !B !A)+(!D !C !B A)+(!D !C B !A)+(!D !C B A)+(!D C !B !A)+(!D C !B A)+(!D C B !A)+(!D C B A)), LSE_LINE_FILE_ID=3, LSE_LCOL=13, LSE_RCOL=44, LSE_LLINE=32, LSE_RLINE=32 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(11[2:53])
    defparam I1.init = 16'b0000000011111111;
    
endmodule
//
// Verilog Description of module inverter_U982
//

module inverter_U982 (\notGate[113]_keep , \notGate[114] ) /* synthesis syn_module_defined=1 */ ;
    input \notGate[113]_keep ;
    output \notGate[114] ;
    
    wire \notGate[113]_keep  /* synthesis alspreserve=1 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(25[15:22])
    
    LUT4 I1 (.A(\notGate[113]_keep ), .B(\notGate[113]_keep ), .C(\notGate[113]_keep ), 
         .D(\notGate[113]_keep ), .Z(\notGate[114] )) /* synthesis syn_instantiated=1, lut_function=((!D !C !B !A)+(!D !C !B A)+(!D !C B !A)+(!D !C B A)+(!D C !B !A)+(!D C !B A)+(!D C B !A)+(!D C B A)), LSE_LINE_FILE_ID=3, LSE_LCOL=13, LSE_RCOL=44, LSE_LLINE=32, LSE_RLINE=32 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(11[2:53])
    defparam I1.init = 16'b0000000011111111;
    
endmodule
//
// Verilog Description of module inverter_U983
//

module inverter_U983 (\notGate[112]_keep , \notGate[113] ) /* synthesis syn_module_defined=1 */ ;
    input \notGate[112]_keep ;
    output \notGate[113] ;
    
    wire \notGate[112]_keep  /* synthesis alspreserve=1 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(25[15:22])
    
    LUT4 I1 (.A(\notGate[112]_keep ), .B(\notGate[112]_keep ), .C(\notGate[112]_keep ), 
         .D(\notGate[112]_keep ), .Z(\notGate[113] )) /* synthesis syn_instantiated=1, lut_function=((!D !C !B !A)+(!D !C !B A)+(!D !C B !A)+(!D !C B A)+(!D C !B !A)+(!D C !B A)+(!D C B !A)+(!D C B A)), LSE_LINE_FILE_ID=3, LSE_LCOL=13, LSE_RCOL=44, LSE_LLINE=32, LSE_RLINE=32 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(11[2:53])
    defparam I1.init = 16'b0000000011111111;
    
endmodule
//
// Verilog Description of module inverter_U984
//

module inverter_U984 (\notGate[111]_keep , \notGate[112] ) /* synthesis syn_module_defined=1 */ ;
    input \notGate[111]_keep ;
    output \notGate[112] ;
    
    wire \notGate[111]_keep  /* synthesis alspreserve=1 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(25[15:22])
    
    LUT4 I1 (.A(\notGate[111]_keep ), .B(\notGate[111]_keep ), .C(\notGate[111]_keep ), 
         .D(\notGate[111]_keep ), .Z(\notGate[112] )) /* synthesis syn_instantiated=1, lut_function=((!D !C !B !A)+(!D !C !B A)+(!D !C B !A)+(!D !C B A)+(!D C !B !A)+(!D C !B A)+(!D C B !A)+(!D C B A)), LSE_LINE_FILE_ID=3, LSE_LCOL=13, LSE_RCOL=44, LSE_LLINE=32, LSE_RLINE=32 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(11[2:53])
    defparam I1.init = 16'b0000000011111111;
    
endmodule
//
// Verilog Description of module inverter_U985
//

module inverter_U985 (\notGate[110]_keep , \notGate[111] ) /* synthesis syn_module_defined=1 */ ;
    input \notGate[110]_keep ;
    output \notGate[111] ;
    
    wire \notGate[110]_keep  /* synthesis alspreserve=1 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(25[15:22])
    
    LUT4 I1 (.A(\notGate[110]_keep ), .B(\notGate[110]_keep ), .C(\notGate[110]_keep ), 
         .D(\notGate[110]_keep ), .Z(\notGate[111] )) /* synthesis syn_instantiated=1, lut_function=((!D !C !B !A)+(!D !C !B A)+(!D !C B !A)+(!D !C B A)+(!D C !B !A)+(!D C !B A)+(!D C B !A)+(!D C B A)), LSE_LINE_FILE_ID=3, LSE_LCOL=13, LSE_RCOL=44, LSE_LLINE=32, LSE_RLINE=32 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(11[2:53])
    defparam I1.init = 16'b0000000011111111;
    
endmodule
//
// Verilog Description of module inverter_U986
//

module inverter_U986 (\notGate[109]_keep , \notGate[110] ) /* synthesis syn_module_defined=1 */ ;
    input \notGate[109]_keep ;
    output \notGate[110] ;
    
    wire \notGate[109]_keep  /* synthesis alspreserve=1 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(25[15:22])
    
    LUT4 I1 (.A(\notGate[109]_keep ), .B(\notGate[109]_keep ), .C(\notGate[109]_keep ), 
         .D(\notGate[109]_keep ), .Z(\notGate[110] )) /* synthesis syn_instantiated=1, lut_function=((!D !C !B !A)+(!D !C !B A)+(!D !C B !A)+(!D !C B A)+(!D C !B !A)+(!D C !B A)+(!D C B !A)+(!D C B A)), LSE_LINE_FILE_ID=3, LSE_LCOL=13, LSE_RCOL=44, LSE_LLINE=32, LSE_RLINE=32 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(11[2:53])
    defparam I1.init = 16'b0000000011111111;
    
endmodule
//
// Verilog Description of module inverter_U987
//

module inverter_U987 (\notGate[9]_keep , \notGate[10] ) /* synthesis syn_module_defined=1 */ ;
    input \notGate[9]_keep ;
    output \notGate[10] ;
    
    wire \notGate[9]_keep  /* synthesis alspreserve=1 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(25[15:22])
    
    LUT4 I1 (.A(\notGate[9]_keep ), .B(\notGate[9]_keep ), .C(\notGate[9]_keep ), 
         .D(\notGate[9]_keep ), .Z(\notGate[10] )) /* synthesis syn_instantiated=1, lut_function=((!D !C !B !A)+(!D !C !B A)+(!D !C B !A)+(!D !C B A)+(!D C !B !A)+(!D C !B A)+(!D C B !A)+(!D C B A)), LSE_LINE_FILE_ID=3, LSE_LCOL=13, LSE_RCOL=44, LSE_LLINE=32, LSE_RLINE=32 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(11[2:53])
    defparam I1.init = 16'b0000000011111111;
    
endmodule
//
// Verilog Description of module inverter_U988
//

module inverter_U988 (\notGate[108]_keep , \notGate[109] ) /* synthesis syn_module_defined=1 */ ;
    input \notGate[108]_keep ;
    output \notGate[109] ;
    
    wire \notGate[108]_keep  /* synthesis alspreserve=1 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(25[15:22])
    
    LUT4 I1 (.A(\notGate[108]_keep ), .B(\notGate[108]_keep ), .C(\notGate[108]_keep ), 
         .D(\notGate[108]_keep ), .Z(\notGate[109] )) /* synthesis syn_instantiated=1, lut_function=((!D !C !B !A)+(!D !C !B A)+(!D !C B !A)+(!D !C B A)+(!D C !B !A)+(!D C !B A)+(!D C B !A)+(!D C B A)), LSE_LINE_FILE_ID=3, LSE_LCOL=13, LSE_RCOL=44, LSE_LLINE=32, LSE_RLINE=32 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(11[2:53])
    defparam I1.init = 16'b0000000011111111;
    
endmodule
//
// Verilog Description of module inverter_U989
//

module inverter_U989 (\notGate[107]_keep , \notGate[108] ) /* synthesis syn_module_defined=1 */ ;
    input \notGate[107]_keep ;
    output \notGate[108] ;
    
    wire \notGate[107]_keep  /* synthesis alspreserve=1 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(25[15:22])
    
    LUT4 I1 (.A(\notGate[107]_keep ), .B(\notGate[107]_keep ), .C(\notGate[107]_keep ), 
         .D(\notGate[107]_keep ), .Z(\notGate[108] )) /* synthesis syn_instantiated=1, lut_function=((!D !C !B !A)+(!D !C !B A)+(!D !C B !A)+(!D !C B A)+(!D C !B !A)+(!D C !B A)+(!D C B !A)+(!D C B A)), LSE_LINE_FILE_ID=3, LSE_LCOL=13, LSE_RCOL=44, LSE_LLINE=32, LSE_RLINE=32 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(11[2:53])
    defparam I1.init = 16'b0000000011111111;
    
endmodule
//
// Verilog Description of module inverter_U990
//

module inverter_U990 (\notGate[106]_keep , \notGate[107] ) /* synthesis syn_module_defined=1 */ ;
    input \notGate[106]_keep ;
    output \notGate[107] ;
    
    wire \notGate[106]_keep  /* synthesis alspreserve=1 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(25[15:22])
    
    LUT4 I1 (.A(\notGate[106]_keep ), .B(\notGate[106]_keep ), .C(\notGate[106]_keep ), 
         .D(\notGate[106]_keep ), .Z(\notGate[107] )) /* synthesis syn_instantiated=1, lut_function=((!D !C !B !A)+(!D !C !B A)+(!D !C B !A)+(!D !C B A)+(!D C !B !A)+(!D C !B A)+(!D C B !A)+(!D C B A)), LSE_LINE_FILE_ID=3, LSE_LCOL=13, LSE_RCOL=44, LSE_LLINE=32, LSE_RLINE=32 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(11[2:53])
    defparam I1.init = 16'b0000000011111111;
    
endmodule
//
// Verilog Description of module inverter_U991
//

module inverter_U991 (\notGate[105]_keep , \notGate[106] ) /* synthesis syn_module_defined=1 */ ;
    input \notGate[105]_keep ;
    output \notGate[106] ;
    
    wire \notGate[105]_keep  /* synthesis alspreserve=1 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(25[15:22])
    
    LUT4 I1 (.A(\notGate[105]_keep ), .B(\notGate[105]_keep ), .C(\notGate[105]_keep ), 
         .D(\notGate[105]_keep ), .Z(\notGate[106] )) /* synthesis syn_instantiated=1, lut_function=((!D !C !B !A)+(!D !C !B A)+(!D !C B !A)+(!D !C B A)+(!D C !B !A)+(!D C !B A)+(!D C B !A)+(!D C B A)), LSE_LINE_FILE_ID=3, LSE_LCOL=13, LSE_RCOL=44, LSE_LLINE=32, LSE_RLINE=32 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(11[2:53])
    defparam I1.init = 16'b0000000011111111;
    
endmodule
//
// Verilog Description of module inverter_U992
//

module inverter_U992 (\notGate[104]_keep , \notGate[105] ) /* synthesis syn_module_defined=1 */ ;
    input \notGate[104]_keep ;
    output \notGate[105] ;
    
    wire \notGate[104]_keep  /* synthesis alspreserve=1 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(25[15:22])
    
    LUT4 I1 (.A(\notGate[104]_keep ), .B(\notGate[104]_keep ), .C(\notGate[104]_keep ), 
         .D(\notGate[104]_keep ), .Z(\notGate[105] )) /* synthesis syn_instantiated=1, lut_function=((!D !C !B !A)+(!D !C !B A)+(!D !C B !A)+(!D !C B A)+(!D C !B !A)+(!D C !B A)+(!D C B !A)+(!D C B A)), LSE_LINE_FILE_ID=3, LSE_LCOL=13, LSE_RCOL=44, LSE_LLINE=32, LSE_RLINE=32 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(11[2:53])
    defparam I1.init = 16'b0000000011111111;
    
endmodule
//
// Verilog Description of module inverter_U993
//

module inverter_U993 (\notGate[103]_keep , \notGate[104] ) /* synthesis syn_module_defined=1 */ ;
    input \notGate[103]_keep ;
    output \notGate[104] ;
    
    wire \notGate[103]_keep  /* synthesis alspreserve=1 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(25[15:22])
    
    LUT4 I1 (.A(\notGate[103]_keep ), .B(\notGate[103]_keep ), .C(\notGate[103]_keep ), 
         .D(\notGate[103]_keep ), .Z(\notGate[104] )) /* synthesis syn_instantiated=1, lut_function=((!D !C !B !A)+(!D !C !B A)+(!D !C B !A)+(!D !C B A)+(!D C !B !A)+(!D C !B A)+(!D C B !A)+(!D C B A)), LSE_LINE_FILE_ID=3, LSE_LCOL=13, LSE_RCOL=44, LSE_LLINE=32, LSE_RLINE=32 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(11[2:53])
    defparam I1.init = 16'b0000000011111111;
    
endmodule
//
// Verilog Description of module inverter_U994
//

module inverter_U994 (\notGate[102]_keep , \notGate[103] ) /* synthesis syn_module_defined=1 */ ;
    input \notGate[102]_keep ;
    output \notGate[103] ;
    
    wire \notGate[102]_keep  /* synthesis alspreserve=1 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(25[15:22])
    
    LUT4 I1 (.A(\notGate[102]_keep ), .B(\notGate[102]_keep ), .C(\notGate[102]_keep ), 
         .D(\notGate[102]_keep ), .Z(\notGate[103] )) /* synthesis syn_instantiated=1, lut_function=((!D !C !B !A)+(!D !C !B A)+(!D !C B !A)+(!D !C B A)+(!D C !B !A)+(!D C !B A)+(!D C B !A)+(!D C B A)), LSE_LINE_FILE_ID=3, LSE_LCOL=13, LSE_RCOL=44, LSE_LLINE=32, LSE_RLINE=32 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(11[2:53])
    defparam I1.init = 16'b0000000011111111;
    
endmodule
//
// Verilog Description of module inverter_U995
//

module inverter_U995 (\notGate[101]_keep , \notGate[102] ) /* synthesis syn_module_defined=1 */ ;
    input \notGate[101]_keep ;
    output \notGate[102] ;
    
    wire \notGate[101]_keep  /* synthesis alspreserve=1 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(25[15:22])
    
    LUT4 I1 (.A(\notGate[101]_keep ), .B(\notGate[101]_keep ), .C(\notGate[101]_keep ), 
         .D(\notGate[101]_keep ), .Z(\notGate[102] )) /* synthesis syn_instantiated=1, lut_function=((!D !C !B !A)+(!D !C !B A)+(!D !C B !A)+(!D !C B A)+(!D C !B !A)+(!D C !B A)+(!D C B !A)+(!D C B A)), LSE_LINE_FILE_ID=3, LSE_LCOL=13, LSE_RCOL=44, LSE_LLINE=32, LSE_RLINE=32 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(11[2:53])
    defparam I1.init = 16'b0000000011111111;
    
endmodule
//
// Verilog Description of module inverter_U996
//

module inverter_U996 (\notGate[100]_keep , \notGate[101] ) /* synthesis syn_module_defined=1 */ ;
    input \notGate[100]_keep ;
    output \notGate[101] ;
    
    wire \notGate[100]_keep  /* synthesis alspreserve=1 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(25[15:22])
    
    LUT4 I1 (.A(\notGate[100]_keep ), .B(\notGate[100]_keep ), .C(\notGate[100]_keep ), 
         .D(\notGate[100]_keep ), .Z(\notGate[101] )) /* synthesis syn_instantiated=1, lut_function=((!D !C !B !A)+(!D !C !B A)+(!D !C B !A)+(!D !C B A)+(!D C !B !A)+(!D C !B A)+(!D C B !A)+(!D C B A)), LSE_LINE_FILE_ID=3, LSE_LCOL=13, LSE_RCOL=44, LSE_LLINE=32, LSE_RLINE=32 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(11[2:53])
    defparam I1.init = 16'b0000000011111111;
    
endmodule
//
// Verilog Description of module inverter_U997
//

module inverter_U997 (\notGate[99]_keep , \notGate[100] ) /* synthesis syn_module_defined=1 */ ;
    input \notGate[99]_keep ;
    output \notGate[100] ;
    
    wire \notGate[99]_keep  /* synthesis alspreserve=1 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(25[15:22])
    
    LUT4 I1 (.A(\notGate[99]_keep ), .B(\notGate[99]_keep ), .C(\notGate[99]_keep ), 
         .D(\notGate[99]_keep ), .Z(\notGate[100] )) /* synthesis syn_instantiated=1, lut_function=((!D !C !B !A)+(!D !C !B A)+(!D !C B !A)+(!D !C B A)+(!D C !B !A)+(!D C !B A)+(!D C B !A)+(!D C B A)), LSE_LINE_FILE_ID=3, LSE_LCOL=13, LSE_RCOL=44, LSE_LLINE=32, LSE_RLINE=32 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(11[2:53])
    defparam I1.init = 16'b0000000011111111;
    
endmodule
//
// Verilog Description of module inverter_U998
//

module inverter_U998 (\notGate[999]_keep , \notGate[1000] ) /* synthesis syn_module_defined=1 */ ;
    input \notGate[999]_keep ;
    output \notGate[1000] ;
    
    wire \notGate[999]_keep  /* synthesis alspreserve=1 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(25[15:22])
    
    LUT4 I1 (.A(\notGate[999]_keep ), .B(\notGate[999]_keep ), .C(\notGate[999]_keep ), 
         .D(\notGate[999]_keep ), .Z(\notGate[1000] )) /* synthesis syn_instantiated=1, lut_function=((!D !C !B !A)+(!D !C !B A)+(!D !C B !A)+(!D !C B A)+(!D C !B !A)+(!D C !B A)+(!D C B !A)+(!D C B A)), LSE_LINE_FILE_ID=3, LSE_LCOL=13, LSE_RCOL=44, LSE_LLINE=32, LSE_RLINE=32 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(11[2:53])
    defparam I1.init = 16'b0000000011111111;
    
endmodule
//
// Verilog Description of module PUR
// module not written out since it is a black-box. 
//

//
// Verilog Description of module \RingOscillatorBase(N=3) 
//

module \RingOscillatorBase(N=3)  (out3_c, run_c_c) /* synthesis syn_module_defined=1 */ ;
    output out3_c;
    input run_c_c;
    
    wire [2:0]notGate_2__N_1 /* synthesis alspreserve=1 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(65[10:14])
    wire notGate_1 /* synthesis alspreserve=1 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(45[14:21])
    wire notGate_0 /* synthesis alspreserve=1 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(45[14:21])
    wire and_1 /* synthesis alspreserve=1 */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(46[6:11])
    
    LUT4 i7_1_lut (.A(notGate_1), .Z(out3_c)) /* synthesis lut_function=(!(A)) */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(54[19:34])
    defparam i7_1_lut.init = 16'h5555;
    LUT4 notGate_0__keep_I_0_1_lut (.A(notGate_0), .Z(notGate_1)) /* synthesis lut_function=(!(A)) */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(54[19:34])
    defparam notGate_0__keep_I_0_1_lut.init = 16'h5555;
    LUT4 en_I_0_2_lut (.A(run_c_c), .B(out3_c), .Z(and_1)) /* synthesis lut_function=(A (B)) */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(51[13:30])
    defparam en_I_0_2_lut.init = 16'h8888;
    LUT4 and_1_keep_I_0_1_lut (.A(and_1), .Z(notGate_0)) /* synthesis lut_function=(!(A)) */ ;   // c:/users/mucar/onedrive/documentos/ufrgs/tcc/lattice 2/osc.v(52[18:24])
    defparam and_1_keep_I_0_1_lut.init = 16'h5555;
    
endmodule
